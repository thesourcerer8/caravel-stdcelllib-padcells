magic
tech sky130A
magscale 1 2
timestamp 1608122862
<< locali >>
rect 27611 55811 27645 55913
rect 44815 43639 44849 43809
rect 8935 24599 8969 24769
rect 12155 23511 12189 23613
rect 9119 22559 9153 22729
rect 9303 22491 9337 22593
rect 8567 21471 8601 21641
rect 8693 18241 9119 18275
rect 8785 18173 9061 18207
rect 9027 18071 9061 18173
rect 23931 17527 23965 17833
rect 27795 15963 27829 16133
rect 34695 15963 34729 16201
rect 12247 8415 12281 8517
<< viali >>
rect 9671 56797 9705 56831
rect 29451 56797 29485 56831
rect 2679 56661 2713 56695
rect 56039 56661 56073 56695
rect 16571 56253 16605 56287
rect 6175 56117 6209 56151
rect 27611 55913 27645 55947
rect 27611 55777 27645 55811
rect 27979 55641 28013 55675
rect 37915 55573 37949 55607
rect 52451 55573 52485 55607
rect 18135 54485 18169 54519
rect 21079 54485 21113 54519
rect 43803 54485 43837 54519
rect 1575 54077 1609 54111
rect 23655 53737 23689 53771
rect 18503 53193 18537 53227
rect 13995 52989 14029 53023
rect 11971 52377 12005 52411
rect 33131 52377 33165 52411
rect 7647 52309 7681 52343
rect 39663 52309 39697 52343
rect 10867 51425 10901 51459
rect 18227 50813 18261 50847
rect 28899 50813 28933 50847
rect 33867 49725 33901 49759
rect 48679 49045 48713 49079
rect 23103 48637 23137 48671
rect 34051 48637 34085 48671
rect 46747 47957 46781 47991
rect 34051 46937 34085 46971
rect 33775 46461 33809 46495
rect 58431 46461 58465 46495
rect 48035 46325 48069 46359
rect 2863 45849 2897 45883
rect 9211 45781 9245 45815
rect 20527 45781 20561 45815
rect 32947 45781 32981 45815
rect 20987 45373 21021 45407
rect 29451 45373 29485 45407
rect 39019 45373 39053 45407
rect 36903 44693 36937 44727
rect 13811 44353 13845 44387
rect 30003 44285 30037 44319
rect 36627 44285 36661 44319
rect 38191 44285 38225 44319
rect 42515 44285 42549 44319
rect 44907 43945 44941 43979
rect 44815 43809 44849 43843
rect 53003 43809 53037 43843
rect 37455 43741 37489 43775
rect 51991 43741 52025 43775
rect 6727 43605 6761 43639
rect 44815 43605 44849 43639
rect 15007 43401 15041 43435
rect 1391 43129 1425 43163
rect 9947 43061 9981 43095
rect 9947 42177 9981 42211
rect 36075 42109 36109 42143
rect 19975 41225 20009 41259
rect 7555 41021 7589 41055
rect 11143 41021 11177 41055
rect 6451 40341 6485 40375
rect 55947 40341 55981 40375
rect 4979 40069 5013 40103
rect 14639 40069 14673 40103
rect 57603 40069 57637 40103
rect 41871 39389 41905 39423
rect 21815 39253 21849 39287
rect 36995 39253 37029 39287
rect 56131 39253 56165 39287
rect 23195 39049 23229 39083
rect 26691 38165 26725 38199
rect 21815 37417 21849 37451
rect 25311 37145 25345 37179
rect 11143 37077 11177 37111
rect 26967 37077 27001 37111
rect 45091 37077 45125 37111
rect 19423 36873 19457 36907
rect 53095 36737 53129 36771
rect 4703 36669 4737 36703
rect 11787 36669 11821 36703
rect 15467 36669 15501 36703
rect 35063 36669 35097 36703
rect 6359 35989 6393 36023
rect 38099 35989 38133 36023
rect 38375 35785 38409 35819
rect 4519 35581 4553 35615
rect 55671 35581 55705 35615
rect 16295 34901 16329 34935
rect 43067 34493 43101 34527
rect 6635 33813 6669 33847
rect 4335 32861 4369 32895
rect 11879 32725 11913 32759
rect 54751 31773 54785 31807
rect 11235 31229 11269 31263
rect 36075 31229 36109 31263
rect 54015 30209 54049 30243
rect 17123 30141 17157 30175
rect 29451 30141 29485 30175
rect 48127 30141 48161 30175
rect 48495 30141 48529 30175
rect 15651 29461 15685 29495
rect 3599 29257 3633 29291
rect 30371 29053 30405 29087
rect 27611 28713 27645 28747
rect 25955 28373 25989 28407
rect 34787 28373 34821 28407
rect 37823 27965 37857 27999
rect 38007 26877 38041 26911
rect 21723 26741 21757 26775
rect 43527 26401 43561 26435
rect 29175 26333 29209 26367
rect 49139 26333 49173 26367
rect 25035 26265 25069 26299
rect 34143 26265 34177 26299
rect 13627 25993 13661 26027
rect 10223 25857 10257 25891
rect 42239 25789 42273 25823
rect 51715 25109 51749 25143
rect 8935 24769 8969 24803
rect 2495 24701 2529 24735
rect 8935 24565 8969 24599
rect 43619 24225 43653 24259
rect 28531 24021 28565 24055
rect 7647 23817 7681 23851
rect 18227 23817 18261 23851
rect 12891 23749 12925 23783
rect 19975 23749 20009 23783
rect 12155 23613 12189 23647
rect 12155 23477 12189 23511
rect 9119 22729 9153 22763
rect 9119 22525 9153 22559
rect 9303 22593 9337 22627
rect 55947 22593 55981 22627
rect 36167 22525 36201 22559
rect 9303 22457 9337 22491
rect 2863 22117 2897 22151
rect 17675 21913 17709 21947
rect 46839 21913 46873 21947
rect 21079 21845 21113 21879
rect 47943 21845 47977 21879
rect 8567 21641 8601 21675
rect 8567 21437 8601 21471
rect 30371 21437 30405 21471
rect 56499 20553 56533 20587
rect 10867 20349 10901 20383
rect 42239 19737 42273 19771
rect 40307 19669 40341 19703
rect 5623 19465 5657 19499
rect 7279 19261 7313 19295
rect 35155 18581 35189 18615
rect 44999 18581 45033 18615
rect 2587 18377 2621 18411
rect 8659 18241 8693 18275
rect 9119 18241 9153 18275
rect 8751 18173 8785 18207
rect 47115 18173 47149 18207
rect 54015 18173 54049 18207
rect 9027 18037 9061 18071
rect 23931 17833 23965 17867
rect 35431 17629 35465 17663
rect 9395 17493 9429 17527
rect 23931 17493 23965 17527
rect 24207 17493 24241 17527
rect 38191 17493 38225 17527
rect 34695 16201 34729 16235
rect 27795 16133 27829 16167
rect 2955 15997 2989 16031
rect 27887 16065 27921 16099
rect 32671 15997 32705 16031
rect 34603 15997 34637 16031
rect 27795 15929 27829 15963
rect 35063 15997 35097 16031
rect 34695 15929 34729 15963
rect 26691 15385 26725 15419
rect 55947 15317 55981 15351
rect 13075 15045 13109 15079
rect 15191 15045 15225 15079
rect 4059 14909 4093 14943
rect 31199 14909 31233 14943
rect 57695 14909 57729 14943
rect 44631 14433 44665 14467
rect 30831 14297 30865 14331
rect 25771 14229 25805 14263
rect 36995 14229 37029 14263
rect 53003 14229 53037 14263
rect 7003 14025 7037 14059
rect 26047 13957 26081 13991
rect 49875 13753 49909 13787
rect 27795 12937 27829 12971
rect 44723 12937 44757 12971
rect 52911 12869 52945 12903
rect 22183 12733 22217 12767
rect 23839 12733 23873 12767
rect 45827 12733 45861 12767
rect 20343 12393 20377 12427
rect 24391 12257 24425 12291
rect 42239 12257 42273 12291
rect 33315 12053 33349 12087
rect 44447 12053 44481 12087
rect 19055 11645 19089 11679
rect 49415 11645 49449 11679
rect 55947 11645 55981 11679
rect 29819 10761 29853 10795
rect 32579 10013 32613 10047
rect 33775 9945 33809 9979
rect 32303 9877 32337 9911
rect 49139 9877 49173 9911
rect 10039 9469 10073 9503
rect 20803 9469 20837 9503
rect 48403 8585 48437 8619
rect 12247 8517 12281 8551
rect 39847 8517 39881 8551
rect 3967 8449 4001 8483
rect 12247 8381 12281 8415
rect 47115 8381 47149 8415
rect 49323 7769 49357 7803
rect 25127 7701 25161 7735
rect 46287 7701 46321 7735
rect 13995 7293 14029 7327
rect 5439 6613 5473 6647
rect 10407 6205 10441 6239
rect 36535 6205 36569 6239
rect 28347 5865 28381 5899
rect 43527 5593 43561 5627
rect 18963 5525 18997 5559
rect 47667 4437 47701 4471
rect 7463 4233 7497 4267
rect 52359 3349 52393 3383
rect 58431 3349 58465 3383
rect 18595 3145 18629 3179
rect 7371 2465 7405 2499
rect 19423 2329 19457 2363
rect 50151 2261 50185 2295
<< metal1 >>
rect 4320 59100 4326 59152
rect 4378 59140 4384 59152
rect 6160 59140 6166 59152
rect 4378 59112 6166 59140
rect 4378 59100 4384 59112
rect 6160 59100 6166 59112
rect 6218 59100 6224 59152
rect 45720 59100 45726 59152
rect 45778 59140 45784 59152
rect 45904 59140 45910 59152
rect 45778 59112 45910 59140
rect 45778 59100 45784 59112
rect 45904 59100 45910 59112
rect 45962 59100 45968 59152
rect 56760 57876 56766 57928
rect 56818 57916 56824 57928
rect 56852 57916 56858 57928
rect 56818 57888 56858 57916
rect 56818 57876 56824 57888
rect 56852 57876 56858 57888
rect 56910 57876 56916 57928
rect 34680 57808 34686 57860
rect 34738 57848 34744 57860
rect 34864 57848 34870 57860
rect 34738 57820 34870 57848
rect 34738 57808 34744 57820
rect 34864 57808 34870 57820
rect 34922 57808 34928 57860
rect 1086 57690 58862 57712
rect 1086 57638 4228 57690
rect 4280 57638 4292 57690
rect 4344 57638 4356 57690
rect 4408 57638 4420 57690
rect 4472 57638 34948 57690
rect 35000 57638 35012 57690
rect 35064 57638 35076 57690
rect 35128 57638 35140 57690
rect 35192 57638 58862 57690
rect 1086 57616 58862 57638
rect 1086 57146 58862 57168
rect 1086 57094 19588 57146
rect 19640 57094 19652 57146
rect 19704 57094 19716 57146
rect 19768 57094 19780 57146
rect 19832 57094 50308 57146
rect 50360 57094 50372 57146
rect 50424 57094 50436 57146
rect 50488 57094 50500 57146
rect 50552 57094 58862 57146
rect 1086 57072 58862 57094
rect 9659 56831 9717 56837
rect 9659 56797 9671 56831
rect 9705 56828 9717 56831
rect 23732 56828 23738 56840
rect 9705 56800 23738 56828
rect 9705 56797 9717 56800
rect 9659 56791 9717 56797
rect 23732 56788 23738 56800
rect 23790 56788 23796 56840
rect 29436 56828 29442 56840
rect 29397 56800 29442 56828
rect 29436 56788 29442 56800
rect 29494 56788 29500 56840
rect 39464 56720 39470 56772
rect 39522 56760 39528 56772
rect 44892 56760 44898 56772
rect 39522 56732 44898 56760
rect 39522 56720 39528 56732
rect 44892 56720 44898 56732
rect 44950 56720 44956 56772
rect 2667 56695 2725 56701
rect 2667 56661 2679 56695
rect 2713 56692 2725 56695
rect 15820 56692 15826 56704
rect 2713 56664 15826 56692
rect 2713 56661 2725 56664
rect 2667 56655 2725 56661
rect 15820 56652 15826 56664
rect 15878 56652 15884 56704
rect 26032 56652 26038 56704
rect 26090 56692 26096 56704
rect 56027 56695 56085 56701
rect 56027 56692 56039 56695
rect 26090 56664 56039 56692
rect 26090 56652 26096 56664
rect 56027 56661 56039 56664
rect 56073 56661 56085 56695
rect 56027 56655 56085 56661
rect 1086 56602 58862 56624
rect 1086 56550 4228 56602
rect 4280 56550 4292 56602
rect 4344 56550 4356 56602
rect 4408 56550 4420 56602
rect 4472 56550 34948 56602
rect 35000 56550 35012 56602
rect 35064 56550 35076 56602
rect 35128 56550 35140 56602
rect 35192 56550 58862 56602
rect 1086 56528 58862 56550
rect 640 56448 646 56500
rect 698 56488 704 56500
rect 1192 56488 1198 56500
rect 698 56460 1198 56488
rect 698 56448 704 56460
rect 1192 56448 1198 56460
rect 1250 56448 1256 56500
rect 1744 56448 1750 56500
rect 1802 56488 1808 56500
rect 2664 56488 2670 56500
rect 1802 56460 2670 56488
rect 1802 56448 1808 56460
rect 2664 56448 2670 56460
rect 2722 56448 2728 56500
rect 13612 56448 13618 56500
rect 13670 56488 13676 56500
rect 13670 56460 21202 56488
rect 13670 56448 13676 56460
rect 180 56380 186 56432
rect 238 56420 244 56432
rect 1284 56420 1290 56432
rect 238 56392 1290 56420
rect 238 56380 244 56392
rect 1284 56380 1290 56392
rect 1342 56380 1348 56432
rect 14440 56380 14446 56432
rect 14498 56420 14504 56432
rect 21064 56420 21070 56432
rect 14498 56392 21070 56420
rect 14498 56380 14504 56392
rect 21064 56380 21070 56392
rect 21122 56380 21128 56432
rect 21174 56420 21202 56460
rect 23732 56448 23738 56500
rect 23790 56488 23796 56500
rect 23790 56460 31874 56488
rect 23790 56448 23796 56460
rect 28056 56420 28062 56432
rect 21174 56392 28062 56420
rect 28056 56380 28062 56392
rect 28114 56380 28120 56432
rect 28148 56380 28154 56432
rect 28206 56420 28212 56432
rect 31184 56420 31190 56432
rect 28206 56392 31190 56420
rect 28206 56380 28212 56392
rect 31184 56380 31190 56392
rect 31242 56380 31248 56432
rect 31846 56420 31874 56460
rect 31920 56448 31926 56500
rect 31978 56488 31984 56500
rect 35968 56488 35974 56500
rect 31978 56460 35974 56488
rect 31978 56448 31984 56460
rect 35968 56448 35974 56460
rect 36026 56448 36032 56500
rect 36060 56448 36066 56500
rect 36118 56488 36124 56500
rect 41396 56488 41402 56500
rect 36118 56460 41402 56488
rect 36118 56448 36124 56460
rect 41396 56448 41402 56460
rect 41454 56448 41460 56500
rect 41488 56448 41494 56500
rect 41546 56488 41552 56500
rect 54828 56488 54834 56500
rect 41546 56460 54834 56488
rect 41546 56448 41552 56460
rect 54828 56448 54834 56460
rect 54886 56448 54892 56500
rect 40108 56420 40114 56432
rect 31846 56392 40114 56420
rect 40108 56380 40114 56392
rect 40166 56380 40172 56432
rect 40200 56380 40206 56432
rect 40258 56420 40264 56432
rect 40258 56392 41258 56420
rect 40258 56380 40264 56392
rect 10852 56312 10858 56364
rect 10910 56352 10916 56364
rect 26676 56352 26682 56364
rect 10910 56324 26682 56352
rect 10910 56312 10916 56324
rect 26676 56312 26682 56324
rect 26734 56312 26740 56364
rect 26768 56312 26774 56364
rect 26826 56352 26832 56364
rect 35876 56352 35882 56364
rect 26826 56324 35882 56352
rect 26826 56312 26832 56324
rect 35876 56312 35882 56324
rect 35934 56312 35940 56364
rect 35968 56312 35974 56364
rect 36026 56352 36032 56364
rect 36026 56324 36198 56352
rect 36026 56312 36032 56324
rect 10576 56244 10582 56296
rect 10634 56284 10640 56296
rect 15912 56284 15918 56296
rect 10634 56256 15918 56284
rect 10634 56244 10640 56256
rect 15912 56244 15918 56256
rect 15970 56244 15976 56296
rect 16559 56287 16617 56293
rect 16559 56253 16571 56287
rect 16605 56284 16617 56287
rect 19960 56284 19966 56296
rect 16605 56256 19966 56284
rect 16605 56253 16617 56256
rect 16559 56247 16617 56253
rect 19960 56244 19966 56256
rect 20018 56244 20024 56296
rect 24008 56244 24014 56296
rect 24066 56284 24072 56296
rect 29436 56284 29442 56296
rect 24066 56256 29442 56284
rect 24066 56244 24072 56256
rect 29436 56244 29442 56256
rect 29494 56244 29500 56296
rect 29712 56244 29718 56296
rect 29770 56284 29776 56296
rect 32932 56284 32938 56296
rect 29770 56256 32938 56284
rect 29770 56244 29776 56256
rect 32932 56244 32938 56256
rect 32990 56244 32996 56296
rect 33024 56244 33030 56296
rect 33082 56284 33088 56296
rect 36060 56284 36066 56296
rect 33082 56256 36066 56284
rect 33082 56244 33088 56256
rect 36060 56244 36066 56256
rect 36118 56244 36124 56296
rect 36170 56284 36198 56324
rect 36520 56312 36526 56364
rect 36578 56352 36584 56364
rect 41120 56352 41126 56364
rect 36578 56324 41126 56352
rect 36578 56312 36584 56324
rect 41120 56312 41126 56324
rect 41178 56312 41184 56364
rect 41230 56352 41258 56392
rect 41304 56380 41310 56432
rect 41362 56420 41368 56432
rect 51148 56420 51154 56432
rect 41362 56392 51154 56420
rect 41362 56380 41368 56392
rect 51148 56380 51154 56392
rect 51206 56380 51212 56432
rect 52712 56352 52718 56364
rect 41230 56324 52718 56352
rect 52712 56312 52718 56324
rect 52770 56312 52776 56364
rect 40660 56284 40666 56296
rect 36170 56256 40666 56284
rect 40660 56244 40666 56256
rect 40718 56244 40724 56296
rect 40752 56244 40758 56296
rect 40810 56284 40816 56296
rect 57496 56284 57502 56296
rect 40810 56256 57502 56284
rect 40810 56244 40816 56256
rect 57496 56244 57502 56256
rect 57554 56244 57560 56296
rect 4044 56176 4050 56228
rect 4102 56216 4108 56228
rect 16464 56216 16470 56228
rect 4102 56188 16470 56216
rect 4102 56176 4108 56188
rect 16464 56176 16470 56188
rect 16522 56176 16528 56228
rect 21616 56176 21622 56228
rect 21674 56216 21680 56228
rect 26860 56216 26866 56228
rect 21674 56188 26866 56216
rect 21674 56176 21680 56188
rect 26860 56176 26866 56188
rect 26918 56176 26924 56228
rect 27044 56176 27050 56228
rect 27102 56216 27108 56228
rect 31552 56216 31558 56228
rect 27102 56188 31558 56216
rect 27102 56176 27108 56188
rect 31552 56176 31558 56188
rect 31610 56176 31616 56228
rect 31644 56176 31650 56228
rect 31702 56216 31708 56228
rect 31702 56188 33162 56216
rect 31702 56176 31708 56188
rect 6163 56151 6221 56157
rect 6163 56117 6175 56151
rect 6209 56148 6221 56151
rect 33024 56148 33030 56160
rect 6209 56120 33030 56148
rect 6209 56117 6221 56120
rect 6163 56111 6221 56117
rect 33024 56108 33030 56120
rect 33082 56108 33088 56160
rect 33134 56148 33162 56188
rect 33208 56176 33214 56228
rect 33266 56216 33272 56228
rect 33266 56188 41534 56216
rect 33266 56176 33272 56188
rect 41396 56148 41402 56160
rect 33134 56120 41402 56148
rect 41396 56108 41402 56120
rect 41454 56108 41460 56160
rect 41506 56148 41534 56188
rect 41580 56176 41586 56228
rect 41638 56216 41644 56228
rect 43236 56216 43242 56228
rect 41638 56188 43242 56216
rect 41638 56176 41644 56188
rect 43236 56176 43242 56188
rect 43294 56176 43300 56228
rect 44156 56176 44162 56228
rect 44214 56216 44220 56228
rect 45352 56216 45358 56228
rect 44214 56188 45358 56216
rect 44214 56176 44220 56188
rect 45352 56176 45358 56188
rect 45410 56176 45416 56228
rect 45444 56176 45450 56228
rect 45502 56216 45508 56228
rect 48572 56216 48578 56228
rect 45502 56188 48578 56216
rect 45502 56176 45508 56188
rect 48572 56176 48578 56188
rect 48630 56176 48636 56228
rect 41672 56148 41678 56160
rect 41506 56120 41678 56148
rect 41672 56108 41678 56120
rect 41730 56108 41736 56160
rect 44892 56108 44898 56160
rect 44950 56148 44956 56160
rect 55932 56148 55938 56160
rect 44950 56120 55938 56148
rect 44950 56108 44956 56120
rect 55932 56108 55938 56120
rect 55990 56108 55996 56160
rect 1086 56058 58862 56080
rect 1086 56006 19588 56058
rect 19640 56006 19652 56058
rect 19704 56006 19716 56058
rect 19768 56006 19780 56058
rect 19832 56006 50308 56058
rect 50360 56006 50372 56058
rect 50424 56006 50436 56058
rect 50488 56006 50500 56058
rect 50552 56006 58862 56058
rect 1086 55984 58862 56006
rect 9840 55904 9846 55956
rect 9898 55944 9904 55956
rect 27599 55947 27657 55953
rect 27599 55944 27611 55947
rect 9898 55916 27611 55944
rect 9898 55904 9904 55916
rect 27599 55913 27611 55916
rect 27645 55913 27657 55947
rect 27599 55907 27657 55913
rect 29804 55904 29810 55956
rect 29862 55944 29868 55956
rect 31644 55944 31650 55956
rect 29862 55916 31650 55944
rect 29862 55904 29868 55916
rect 31644 55904 31650 55916
rect 31702 55904 31708 55956
rect 31736 55904 31742 55956
rect 31794 55944 31800 55956
rect 33208 55944 33214 55956
rect 31794 55916 33214 55944
rect 31794 55904 31800 55916
rect 33208 55904 33214 55916
rect 33266 55904 33272 55956
rect 35416 55904 35422 55956
rect 35474 55944 35480 55956
rect 38636 55944 38642 55956
rect 35474 55916 38642 55944
rect 35474 55904 35480 55916
rect 38636 55904 38642 55916
rect 38694 55904 38700 55956
rect 39648 55904 39654 55956
rect 39706 55944 39712 55956
rect 58048 55944 58054 55956
rect 39706 55916 58054 55944
rect 39706 55904 39712 55916
rect 58048 55904 58054 55916
rect 58106 55904 58112 55956
rect 8092 55836 8098 55888
rect 8150 55876 8156 55888
rect 44156 55876 44162 55888
rect 8150 55848 44162 55876
rect 8150 55836 8156 55848
rect 44156 55836 44162 55848
rect 44214 55836 44220 55888
rect 44708 55836 44714 55888
rect 44766 55876 44772 55888
rect 59060 55876 59066 55888
rect 44766 55848 59066 55876
rect 44766 55836 44772 55848
rect 59060 55836 59066 55848
rect 59118 55836 59124 55888
rect 8552 55768 8558 55820
rect 8610 55808 8616 55820
rect 13060 55808 13066 55820
rect 8610 55780 13066 55808
rect 8610 55768 8616 55780
rect 13060 55768 13066 55780
rect 13118 55768 13124 55820
rect 20144 55768 20150 55820
rect 20202 55808 20208 55820
rect 26216 55808 26222 55820
rect 20202 55780 26222 55808
rect 20202 55768 20208 55780
rect 26216 55768 26222 55780
rect 26274 55768 26280 55820
rect 27599 55811 27657 55817
rect 27599 55777 27611 55811
rect 27645 55808 27657 55811
rect 37532 55808 37538 55820
rect 27645 55780 37538 55808
rect 27645 55777 27657 55780
rect 27599 55771 27657 55777
rect 37532 55768 37538 55780
rect 37590 55768 37596 55820
rect 37624 55768 37630 55820
rect 37682 55808 37688 55820
rect 40568 55808 40574 55820
rect 37682 55780 40574 55808
rect 37682 55768 37688 55780
rect 40568 55768 40574 55780
rect 40626 55768 40632 55820
rect 40660 55768 40666 55820
rect 40718 55808 40724 55820
rect 59612 55808 59618 55820
rect 40718 55780 59618 55808
rect 40718 55768 40724 55780
rect 59612 55768 59618 55780
rect 59670 55768 59676 55820
rect 7264 55700 7270 55752
rect 7322 55740 7328 55752
rect 18028 55740 18034 55752
rect 7322 55712 18034 55740
rect 7322 55700 7328 55712
rect 18028 55700 18034 55712
rect 18086 55700 18092 55752
rect 19408 55700 19414 55752
rect 19466 55740 19472 55752
rect 26768 55740 26774 55752
rect 19466 55712 26774 55740
rect 19466 55700 19472 55712
rect 26768 55700 26774 55712
rect 26826 55700 26832 55752
rect 26860 55700 26866 55752
rect 26918 55740 26924 55752
rect 33852 55740 33858 55752
rect 26918 55712 33858 55740
rect 26918 55700 26924 55712
rect 33852 55700 33858 55712
rect 33910 55700 33916 55752
rect 33944 55700 33950 55752
rect 34002 55740 34008 55752
rect 34002 55712 35462 55740
rect 34002 55700 34008 55712
rect 10484 55632 10490 55684
rect 10542 55672 10548 55684
rect 17476 55672 17482 55684
rect 10542 55644 17482 55672
rect 10542 55632 10548 55644
rect 17476 55632 17482 55644
rect 17534 55632 17540 55684
rect 18672 55632 18678 55684
rect 18730 55672 18736 55684
rect 22720 55672 22726 55684
rect 18730 55644 22726 55672
rect 18730 55632 18736 55644
rect 22720 55632 22726 55644
rect 22778 55632 22784 55684
rect 26216 55632 26222 55684
rect 26274 55672 26280 55684
rect 27504 55672 27510 55684
rect 26274 55644 27510 55672
rect 26274 55632 26280 55644
rect 27504 55632 27510 55644
rect 27562 55632 27568 55684
rect 27967 55675 28025 55681
rect 27967 55641 27979 55675
rect 28013 55672 28025 55675
rect 31920 55672 31926 55684
rect 28013 55644 31926 55672
rect 28013 55641 28025 55644
rect 27967 55635 28025 55641
rect 31920 55632 31926 55644
rect 31978 55632 31984 55684
rect 32012 55632 32018 55684
rect 32070 55672 32076 55684
rect 35324 55672 35330 55684
rect 32070 55644 35330 55672
rect 32070 55632 32076 55644
rect 35324 55632 35330 55644
rect 35382 55632 35388 55684
rect 35434 55672 35462 55712
rect 35876 55700 35882 55752
rect 35934 55740 35940 55752
rect 38544 55740 38550 55752
rect 35934 55712 38550 55740
rect 35934 55700 35940 55712
rect 38544 55700 38550 55712
rect 38602 55700 38608 55752
rect 38636 55700 38642 55752
rect 38694 55740 38700 55752
rect 53264 55740 53270 55752
rect 38694 55712 53270 55740
rect 38694 55700 38700 55712
rect 53264 55700 53270 55712
rect 53322 55700 53328 55752
rect 37072 55672 37078 55684
rect 35434 55644 37078 55672
rect 37072 55632 37078 55644
rect 37130 55632 37136 55684
rect 38084 55632 38090 55684
rect 38142 55672 38148 55684
rect 42224 55672 42230 55684
rect 38142 55644 42230 55672
rect 38142 55632 38148 55644
rect 42224 55632 42230 55644
rect 42282 55632 42288 55684
rect 44616 55632 44622 55684
rect 44674 55672 44680 55684
rect 54368 55672 54374 55684
rect 44674 55644 54374 55672
rect 44674 55632 44680 55644
rect 54368 55632 54374 55644
rect 54426 55632 54432 55684
rect 13244 55564 13250 55616
rect 13302 55604 13308 55616
rect 20972 55604 20978 55616
rect 13302 55576 20978 55604
rect 13302 55564 13308 55576
rect 20972 55564 20978 55576
rect 21030 55564 21036 55616
rect 21064 55564 21070 55616
rect 21122 55604 21128 55616
rect 23272 55604 23278 55616
rect 21122 55576 23278 55604
rect 21122 55564 21128 55576
rect 23272 55564 23278 55576
rect 23330 55564 23336 55616
rect 25940 55564 25946 55616
rect 25998 55604 26004 55616
rect 27412 55604 27418 55616
rect 25998 55576 27418 55604
rect 25998 55564 26004 55576
rect 27412 55564 27418 55576
rect 27470 55564 27476 55616
rect 27596 55564 27602 55616
rect 27654 55604 27660 55616
rect 31092 55604 31098 55616
rect 27654 55576 31098 55604
rect 27654 55564 27660 55576
rect 31092 55564 31098 55576
rect 31150 55564 31156 55616
rect 31184 55564 31190 55616
rect 31242 55604 31248 55616
rect 37903 55607 37961 55613
rect 37903 55604 37915 55607
rect 31242 55576 37915 55604
rect 31242 55564 31248 55576
rect 37903 55573 37915 55576
rect 37949 55573 37961 55607
rect 37903 55567 37961 55573
rect 38268 55564 38274 55616
rect 38326 55604 38332 55616
rect 41396 55604 41402 55616
rect 38326 55576 41402 55604
rect 38326 55564 38332 55576
rect 41396 55564 41402 55576
rect 41454 55564 41460 55616
rect 41488 55564 41494 55616
rect 41546 55604 41552 55616
rect 47008 55604 47014 55616
rect 41546 55576 47014 55604
rect 41546 55564 41552 55576
rect 47008 55564 47014 55576
rect 47066 55564 47072 55616
rect 52436 55604 52442 55616
rect 52397 55576 52442 55604
rect 52436 55564 52442 55576
rect 52494 55564 52500 55616
rect 1086 55514 58862 55536
rect 1086 55462 4228 55514
rect 4280 55462 4292 55514
rect 4344 55462 4356 55514
rect 4408 55462 4420 55514
rect 4472 55462 34948 55514
rect 35000 55462 35012 55514
rect 35064 55462 35076 55514
rect 35128 55462 35140 55514
rect 35192 55462 58862 55514
rect 1086 55440 58862 55462
rect 17568 55360 17574 55412
rect 17626 55400 17632 55412
rect 20696 55400 20702 55412
rect 17626 55372 20702 55400
rect 17626 55360 17632 55372
rect 20696 55360 20702 55372
rect 20754 55360 20760 55412
rect 23364 55360 23370 55412
rect 23422 55400 23428 55412
rect 30908 55400 30914 55412
rect 23422 55372 30914 55400
rect 23422 55360 23428 55372
rect 30908 55360 30914 55372
rect 30966 55360 30972 55412
rect 31460 55400 31466 55412
rect 31018 55372 31466 55400
rect 4872 55292 4878 55344
rect 4930 55332 4936 55344
rect 6252 55332 6258 55344
rect 4930 55304 6258 55332
rect 4930 55292 4936 55304
rect 6252 55292 6258 55304
rect 6310 55292 6316 55344
rect 6436 55292 6442 55344
rect 6494 55332 6500 55344
rect 8184 55332 8190 55344
rect 6494 55304 8190 55332
rect 6494 55292 6500 55304
rect 8184 55292 8190 55304
rect 8242 55292 8248 55344
rect 14992 55292 14998 55344
rect 15050 55332 15056 55344
rect 17016 55332 17022 55344
rect 15050 55304 17022 55332
rect 15050 55292 15056 55304
rect 17016 55292 17022 55304
rect 17074 55292 17080 55344
rect 20052 55292 20058 55344
rect 20110 55332 20116 55344
rect 20110 55304 20742 55332
rect 20110 55292 20116 55304
rect 2756 55224 2762 55276
rect 2814 55264 2820 55276
rect 3952 55264 3958 55276
rect 2814 55236 3958 55264
rect 2814 55224 2820 55236
rect 3952 55224 3958 55236
rect 4010 55224 4016 55276
rect 5884 55224 5890 55276
rect 5942 55264 5948 55276
rect 6804 55264 6810 55276
rect 5942 55236 6810 55264
rect 5942 55224 5948 55236
rect 6804 55224 6810 55236
rect 6862 55224 6868 55276
rect 6988 55224 6994 55276
rect 7046 55264 7052 55276
rect 8000 55264 8006 55276
rect 7046 55236 8006 55264
rect 7046 55224 7052 55236
rect 8000 55224 8006 55236
rect 8058 55224 8064 55276
rect 8276 55224 8282 55276
rect 8334 55264 8340 55276
rect 9564 55264 9570 55276
rect 8334 55236 9570 55264
rect 8334 55224 8340 55236
rect 9564 55224 9570 55236
rect 9622 55224 9628 55276
rect 11680 55224 11686 55276
rect 11738 55264 11744 55276
rect 12140 55264 12146 55276
rect 11738 55236 12146 55264
rect 11738 55224 11744 55236
rect 12140 55224 12146 55236
rect 12198 55224 12204 55276
rect 13796 55224 13802 55276
rect 13854 55264 13860 55276
rect 15084 55264 15090 55276
rect 13854 55236 15090 55264
rect 13854 55224 13860 55236
rect 15084 55224 15090 55236
rect 15142 55224 15148 55276
rect 18580 55224 18586 55276
rect 18638 55264 18644 55276
rect 19132 55264 19138 55276
rect 18638 55236 19138 55264
rect 18638 55224 18644 55236
rect 19132 55224 19138 55236
rect 19190 55224 19196 55276
rect 19868 55224 19874 55276
rect 19926 55264 19932 55276
rect 20604 55264 20610 55276
rect 19926 55236 20610 55264
rect 19926 55224 19932 55236
rect 20604 55224 20610 55236
rect 20662 55224 20668 55276
rect 20714 55264 20742 55304
rect 20972 55292 20978 55344
rect 21030 55332 21036 55344
rect 24008 55332 24014 55344
rect 21030 55304 24014 55332
rect 21030 55292 21036 55304
rect 24008 55292 24014 55304
rect 24066 55292 24072 55344
rect 29068 55292 29074 55344
rect 29126 55332 29132 55344
rect 30264 55332 30270 55344
rect 29126 55304 30270 55332
rect 29126 55292 29132 55304
rect 30264 55292 30270 55304
rect 30322 55292 30328 55344
rect 20714 55236 24790 55264
rect 24762 55196 24790 55236
rect 24836 55224 24842 55276
rect 24894 55264 24900 55276
rect 26032 55264 26038 55276
rect 24894 55236 26038 55264
rect 24894 55224 24900 55236
rect 26032 55224 26038 55236
rect 26090 55224 26096 55276
rect 26142 55236 28194 55264
rect 26142 55196 26170 55236
rect 24762 55168 26170 55196
rect 28166 55196 28194 55236
rect 28240 55224 28246 55276
rect 28298 55264 28304 55276
rect 29620 55264 29626 55276
rect 28298 55236 29626 55264
rect 28298 55224 28304 55236
rect 29620 55224 29626 55236
rect 29678 55224 29684 55276
rect 31018 55264 31046 55372
rect 31460 55360 31466 55372
rect 31518 55360 31524 55412
rect 31828 55360 31834 55412
rect 31886 55400 31892 55412
rect 31886 55372 32886 55400
rect 31886 55360 31892 55372
rect 31092 55292 31098 55344
rect 31150 55332 31156 55344
rect 32012 55332 32018 55344
rect 31150 55304 32018 55332
rect 31150 55292 31156 55304
rect 32012 55292 32018 55304
rect 32070 55292 32076 55344
rect 32748 55332 32754 55344
rect 32122 55304 32754 55332
rect 32122 55264 32150 55304
rect 32748 55292 32754 55304
rect 32806 55292 32812 55344
rect 32858 55332 32886 55372
rect 32932 55360 32938 55412
rect 32990 55400 32996 55412
rect 36980 55400 36986 55412
rect 32990 55372 36986 55400
rect 32990 55360 32996 55372
rect 36980 55360 36986 55372
rect 37038 55360 37044 55412
rect 37072 55360 37078 55412
rect 37130 55400 37136 55412
rect 41304 55400 41310 55412
rect 37130 55372 41310 55400
rect 37130 55360 37136 55372
rect 41304 55360 41310 55372
rect 41362 55360 41368 55412
rect 41672 55360 41678 55412
rect 41730 55400 41736 55412
rect 43788 55400 43794 55412
rect 41730 55372 43794 55400
rect 41730 55360 41736 55372
rect 43788 55360 43794 55372
rect 43846 55360 43852 55412
rect 43880 55360 43886 55412
rect 43938 55400 43944 55412
rect 46456 55400 46462 55412
rect 43938 55372 46462 55400
rect 43938 55360 43944 55372
rect 46456 55360 46462 55372
rect 46514 55360 46520 55412
rect 39464 55332 39470 55344
rect 32858 55304 39470 55332
rect 39464 55292 39470 55304
rect 39522 55292 39528 55344
rect 43604 55292 43610 55344
rect 43662 55332 43668 55344
rect 50136 55332 50142 55344
rect 43662 55304 50142 55332
rect 43662 55292 43668 55304
rect 50136 55292 50142 55304
rect 50194 55292 50200 55344
rect 29730 55236 31046 55264
rect 31202 55236 32150 55264
rect 29730 55196 29758 55236
rect 28166 55168 29758 55196
rect 31000 55156 31006 55208
rect 31058 55196 31064 55208
rect 31202 55196 31230 55236
rect 32196 55224 32202 55276
rect 32254 55264 32260 55276
rect 33024 55264 33030 55276
rect 32254 55236 33030 55264
rect 32254 55224 32260 55236
rect 33024 55224 33030 55236
rect 33082 55224 33088 55276
rect 33944 55264 33950 55276
rect 33134 55236 33950 55264
rect 31058 55168 31230 55196
rect 31058 55156 31064 55168
rect 32380 55156 32386 55208
rect 32438 55196 32444 55208
rect 33134 55196 33162 55236
rect 33944 55224 33950 55236
rect 34002 55224 34008 55276
rect 34054 55236 35278 55264
rect 32438 55168 33162 55196
rect 32438 55156 32444 55168
rect 33208 55156 33214 55208
rect 33266 55196 33272 55208
rect 34054 55196 34082 55236
rect 33266 55168 34082 55196
rect 33266 55156 33272 55168
rect 30908 55088 30914 55140
rect 30966 55128 30972 55140
rect 32932 55128 32938 55140
rect 30966 55100 32938 55128
rect 30966 55088 30972 55100
rect 32932 55088 32938 55100
rect 32990 55088 32996 55140
rect 35250 55128 35278 55236
rect 35324 55224 35330 55276
rect 35382 55264 35388 55276
rect 41304 55264 41310 55276
rect 35382 55236 41310 55264
rect 35382 55224 35388 55236
rect 41304 55224 41310 55236
rect 41362 55224 41368 55276
rect 41488 55224 41494 55276
rect 41546 55264 41552 55276
rect 51700 55264 51706 55276
rect 41546 55236 51706 55264
rect 41546 55224 41552 55236
rect 51700 55224 51706 55236
rect 51758 55224 51764 55276
rect 43880 55128 43886 55140
rect 35250 55100 43886 55128
rect 43880 55088 43886 55100
rect 43938 55088 43944 55140
rect 33852 55020 33858 55072
rect 33910 55060 33916 55072
rect 37624 55060 37630 55072
rect 33910 55032 37630 55060
rect 33910 55020 33916 55032
rect 37624 55020 37630 55032
rect 37682 55020 37688 55072
rect 1086 54970 58862 54992
rect 1086 54918 19588 54970
rect 19640 54918 19652 54970
rect 19704 54918 19716 54970
rect 19768 54918 19780 54970
rect 19832 54918 50308 54970
rect 50360 54918 50372 54970
rect 50424 54918 50436 54970
rect 50488 54918 50500 54970
rect 50552 54918 58862 54970
rect 1086 54896 58862 54918
rect 19316 54584 19322 54596
rect 11422 54556 19322 54584
rect 4044 54476 4050 54528
rect 4102 54516 4108 54528
rect 11422 54516 11450 54556
rect 19316 54544 19322 54556
rect 19374 54544 19380 54596
rect 18120 54516 18126 54528
rect 4102 54488 11450 54516
rect 18081 54488 18126 54516
rect 4102 54476 4108 54488
rect 18120 54476 18126 54488
rect 18178 54476 18184 54528
rect 21067 54519 21125 54525
rect 21067 54485 21079 54519
rect 21113 54516 21125 54519
rect 22536 54516 22542 54528
rect 21113 54488 22542 54516
rect 21113 54485 21125 54488
rect 21067 54479 21125 54485
rect 22536 54476 22542 54488
rect 22594 54476 22600 54528
rect 23548 54476 23554 54528
rect 23606 54516 23612 54528
rect 43791 54519 43849 54525
rect 43791 54516 43803 54519
rect 23606 54488 43803 54516
rect 23606 54476 23612 54488
rect 43791 54485 43803 54488
rect 43837 54485 43849 54519
rect 43791 54479 43849 54485
rect 1086 54426 58862 54448
rect 1086 54374 4228 54426
rect 4280 54374 4292 54426
rect 4344 54374 4356 54426
rect 4408 54374 4420 54426
rect 4472 54374 34948 54426
rect 35000 54374 35012 54426
rect 35064 54374 35076 54426
rect 35128 54374 35140 54426
rect 35192 54374 58862 54426
rect 1086 54352 58862 54374
rect 22536 54272 22542 54324
rect 22594 54312 22600 54324
rect 48940 54312 48946 54324
rect 22594 54284 48946 54312
rect 22594 54272 22600 54284
rect 48940 54272 48946 54284
rect 48998 54272 49004 54324
rect 21708 54204 21714 54256
rect 21766 54244 21772 54256
rect 27136 54244 27142 54256
rect 21766 54216 27142 54244
rect 21766 54204 21772 54216
rect 27136 54204 27142 54216
rect 27194 54204 27200 54256
rect 1563 54111 1621 54117
rect 1563 54077 1575 54111
rect 1609 54108 1621 54111
rect 22720 54108 22726 54120
rect 1609 54080 22726 54108
rect 1609 54077 1621 54080
rect 1563 54071 1621 54077
rect 22720 54068 22726 54080
rect 22778 54068 22784 54120
rect 1086 53882 58862 53904
rect 1086 53830 19588 53882
rect 19640 53830 19652 53882
rect 19704 53830 19716 53882
rect 19768 53830 19780 53882
rect 19832 53830 50308 53882
rect 50360 53830 50372 53882
rect 50424 53830 50436 53882
rect 50488 53830 50500 53882
rect 50552 53830 58862 53882
rect 1086 53808 58862 53830
rect 23643 53771 23701 53777
rect 23643 53737 23655 53771
rect 23689 53768 23701 53771
rect 30632 53768 30638 53780
rect 23689 53740 30638 53768
rect 23689 53737 23701 53740
rect 23643 53731 23701 53737
rect 30632 53728 30638 53740
rect 30690 53728 30696 53780
rect 1086 53338 58862 53360
rect 1086 53286 4228 53338
rect 4280 53286 4292 53338
rect 4344 53286 4356 53338
rect 4408 53286 4420 53338
rect 4472 53286 34948 53338
rect 35000 53286 35012 53338
rect 35064 53286 35076 53338
rect 35128 53286 35140 53338
rect 35192 53286 58862 53338
rect 1086 53264 58862 53286
rect 18491 53227 18549 53233
rect 18491 53193 18503 53227
rect 18537 53224 18549 53227
rect 23364 53224 23370 53236
rect 18537 53196 23370 53224
rect 18537 53193 18549 53196
rect 18491 53187 18549 53193
rect 23364 53184 23370 53196
rect 23422 53184 23428 53236
rect 39004 53048 39010 53100
rect 39062 53088 39068 53100
rect 39556 53088 39562 53100
rect 39062 53060 39562 53088
rect 39062 53048 39068 53060
rect 39556 53048 39562 53060
rect 39614 53048 39620 53100
rect 12324 52980 12330 53032
rect 12382 53020 12388 53032
rect 13983 53023 14041 53029
rect 13983 53020 13995 53023
rect 12382 52992 13995 53020
rect 12382 52980 12388 52992
rect 13983 52989 13995 52992
rect 14029 52989 14041 53023
rect 13983 52983 14041 52989
rect 1086 52794 58862 52816
rect 1086 52742 19588 52794
rect 19640 52742 19652 52794
rect 19704 52742 19716 52794
rect 19768 52742 19780 52794
rect 19832 52742 50308 52794
rect 50360 52742 50372 52794
rect 50424 52742 50436 52794
rect 50488 52742 50500 52794
rect 50552 52742 58862 52794
rect 1086 52720 58862 52742
rect 5056 52368 5062 52420
rect 5114 52408 5120 52420
rect 11959 52411 12017 52417
rect 11959 52408 11971 52411
rect 5114 52380 11971 52408
rect 5114 52368 5120 52380
rect 11959 52377 11971 52380
rect 12005 52377 12017 52411
rect 11959 52371 12017 52377
rect 33119 52411 33177 52417
rect 33119 52377 33131 52411
rect 33165 52408 33177 52411
rect 35876 52408 35882 52420
rect 33165 52380 35882 52408
rect 33165 52377 33177 52380
rect 33119 52371 33177 52377
rect 35876 52368 35882 52380
rect 35934 52368 35940 52420
rect 7632 52340 7638 52352
rect 7593 52312 7638 52340
rect 7632 52300 7638 52312
rect 7690 52300 7696 52352
rect 39648 52340 39654 52352
rect 39609 52312 39654 52340
rect 39648 52300 39654 52312
rect 39706 52300 39712 52352
rect 1086 52250 58862 52272
rect 1086 52198 4228 52250
rect 4280 52198 4292 52250
rect 4344 52198 4356 52250
rect 4408 52198 4420 52250
rect 4472 52198 34948 52250
rect 35000 52198 35012 52250
rect 35064 52198 35076 52250
rect 35128 52198 35140 52250
rect 35192 52198 58862 52250
rect 1086 52176 58862 52198
rect 1086 51706 58862 51728
rect 1086 51654 19588 51706
rect 19640 51654 19652 51706
rect 19704 51654 19716 51706
rect 19768 51654 19780 51706
rect 19832 51654 50308 51706
rect 50360 51654 50372 51706
rect 50424 51654 50436 51706
rect 50488 51654 50500 51706
rect 50552 51654 58862 51706
rect 1086 51632 58862 51654
rect 10852 51456 10858 51468
rect 10813 51428 10858 51456
rect 10852 51416 10858 51428
rect 10910 51416 10916 51468
rect 1086 51162 58862 51184
rect 1086 51110 4228 51162
rect 4280 51110 4292 51162
rect 4344 51110 4356 51162
rect 4408 51110 4420 51162
rect 4472 51110 34948 51162
rect 35000 51110 35012 51162
rect 35064 51110 35076 51162
rect 35128 51110 35140 51162
rect 35192 51110 58862 51162
rect 1086 51088 58862 51110
rect 13796 51008 13802 51060
rect 13854 51048 13860 51060
rect 14900 51048 14906 51060
rect 13854 51020 14906 51048
rect 13854 51008 13860 51020
rect 14900 51008 14906 51020
rect 14958 51008 14964 51060
rect 18212 50844 18218 50856
rect 18173 50816 18218 50844
rect 18212 50804 18218 50816
rect 18270 50804 18276 50856
rect 28884 50844 28890 50856
rect 28845 50816 28890 50844
rect 28884 50804 28890 50816
rect 28942 50804 28948 50856
rect 1086 50618 58862 50640
rect 1086 50566 19588 50618
rect 19640 50566 19652 50618
rect 19704 50566 19716 50618
rect 19768 50566 19780 50618
rect 19832 50566 50308 50618
rect 50360 50566 50372 50618
rect 50424 50566 50436 50618
rect 50488 50566 50500 50618
rect 50552 50566 58862 50618
rect 1086 50544 58862 50566
rect 1086 50074 58862 50096
rect 1086 50022 4228 50074
rect 4280 50022 4292 50074
rect 4344 50022 4356 50074
rect 4408 50022 4420 50074
rect 4472 50022 34948 50074
rect 35000 50022 35012 50074
rect 35064 50022 35076 50074
rect 35128 50022 35140 50074
rect 35192 50022 58862 50074
rect 1086 50000 58862 50022
rect 16464 49716 16470 49768
rect 16522 49756 16528 49768
rect 33855 49759 33913 49765
rect 33855 49756 33867 49759
rect 16522 49728 33867 49756
rect 16522 49716 16528 49728
rect 33855 49725 33867 49728
rect 33901 49725 33913 49759
rect 33855 49719 33913 49725
rect 1086 49530 58862 49552
rect 1086 49478 19588 49530
rect 19640 49478 19652 49530
rect 19704 49478 19716 49530
rect 19768 49478 19780 49530
rect 19832 49478 50308 49530
rect 50360 49478 50372 49530
rect 50424 49478 50436 49530
rect 50488 49478 50500 49530
rect 50552 49478 58862 49530
rect 1086 49456 58862 49478
rect 18856 49036 18862 49088
rect 18914 49076 18920 49088
rect 48667 49079 48725 49085
rect 48667 49076 48679 49079
rect 18914 49048 48679 49076
rect 18914 49036 18920 49048
rect 48667 49045 48679 49048
rect 48713 49045 48725 49079
rect 48667 49039 48725 49045
rect 1086 48986 58862 49008
rect 1086 48934 4228 48986
rect 4280 48934 4292 48986
rect 4344 48934 4356 48986
rect 4408 48934 4420 48986
rect 4472 48934 34948 48986
rect 35000 48934 35012 48986
rect 35064 48934 35076 48986
rect 35128 48934 35140 48986
rect 35192 48934 58862 48986
rect 1086 48912 58862 48934
rect 13704 48628 13710 48680
rect 13762 48668 13768 48680
rect 23091 48671 23149 48677
rect 23091 48668 23103 48671
rect 13762 48640 23103 48668
rect 13762 48628 13768 48640
rect 23091 48637 23103 48640
rect 23137 48637 23149 48671
rect 34036 48668 34042 48680
rect 33997 48640 34042 48668
rect 23091 48631 23149 48637
rect 34036 48628 34042 48640
rect 34094 48628 34100 48680
rect 1086 48442 58862 48464
rect 1086 48390 19588 48442
rect 19640 48390 19652 48442
rect 19704 48390 19716 48442
rect 19768 48390 19780 48442
rect 19832 48390 50308 48442
rect 50360 48390 50372 48442
rect 50424 48390 50436 48442
rect 50488 48390 50500 48442
rect 50552 48390 58862 48442
rect 1086 48368 58862 48390
rect 8644 48288 8650 48340
rect 8702 48328 8708 48340
rect 8736 48328 8742 48340
rect 8702 48300 8742 48328
rect 8702 48288 8708 48300
rect 8736 48288 8742 48300
rect 8794 48288 8800 48340
rect 18856 48288 18862 48340
rect 18914 48328 18920 48340
rect 18948 48328 18954 48340
rect 18914 48300 18954 48328
rect 18914 48288 18920 48300
rect 18948 48288 18954 48300
rect 19006 48288 19012 48340
rect 24192 48288 24198 48340
rect 24250 48328 24256 48340
rect 26400 48328 26406 48340
rect 24250 48300 26406 48328
rect 24250 48288 24256 48300
rect 26400 48288 26406 48300
rect 26458 48288 26464 48340
rect 29344 48288 29350 48340
rect 29402 48328 29408 48340
rect 30172 48328 30178 48340
rect 29402 48300 30178 48328
rect 29402 48288 29408 48300
rect 30172 48288 30178 48300
rect 30230 48288 30236 48340
rect 34588 48288 34594 48340
rect 34646 48328 34652 48340
rect 34680 48328 34686 48340
rect 34646 48300 34686 48328
rect 34646 48288 34652 48300
rect 34680 48288 34686 48300
rect 34738 48288 34744 48340
rect 37992 48288 37998 48340
rect 38050 48328 38056 48340
rect 38084 48328 38090 48340
rect 38050 48300 38090 48328
rect 38050 48288 38056 48300
rect 38084 48288 38090 48300
rect 38142 48288 38148 48340
rect 35416 48220 35422 48272
rect 35474 48220 35480 48272
rect 51148 48220 51154 48272
rect 51206 48260 51212 48272
rect 51240 48260 51246 48272
rect 51206 48232 51246 48260
rect 51206 48220 51212 48232
rect 51240 48220 51246 48232
rect 51298 48220 51304 48272
rect 35434 48192 35462 48220
rect 35508 48192 35514 48204
rect 35434 48164 35514 48192
rect 35508 48152 35514 48164
rect 35566 48152 35572 48204
rect 34404 47948 34410 48000
rect 34462 47988 34468 48000
rect 46735 47991 46793 47997
rect 46735 47988 46747 47991
rect 34462 47960 46747 47988
rect 34462 47948 34468 47960
rect 46735 47957 46747 47960
rect 46781 47957 46793 47991
rect 46735 47951 46793 47957
rect 1086 47898 58862 47920
rect 1086 47846 4228 47898
rect 4280 47846 4292 47898
rect 4344 47846 4356 47898
rect 4408 47846 4420 47898
rect 4472 47846 34948 47898
rect 35000 47846 35012 47898
rect 35064 47846 35076 47898
rect 35128 47846 35140 47898
rect 35192 47846 58862 47898
rect 1086 47824 58862 47846
rect 1086 47354 58862 47376
rect 1086 47302 19588 47354
rect 19640 47302 19652 47354
rect 19704 47302 19716 47354
rect 19768 47302 19780 47354
rect 19832 47302 50308 47354
rect 50360 47302 50372 47354
rect 50424 47302 50436 47354
rect 50488 47302 50500 47354
rect 50552 47302 58862 47354
rect 1086 47280 58862 47302
rect 26860 47036 26866 47048
rect 26602 47008 26866 47036
rect 26602 46980 26630 47008
rect 26860 46996 26866 47008
rect 26918 46996 26924 47048
rect 10300 46928 10306 46980
rect 10358 46968 10364 46980
rect 10576 46968 10582 46980
rect 10358 46940 10582 46968
rect 10358 46928 10364 46940
rect 10576 46928 10582 46940
rect 10634 46928 10640 46980
rect 17200 46928 17206 46980
rect 17258 46968 17264 46980
rect 17568 46968 17574 46980
rect 17258 46940 17574 46968
rect 17258 46928 17264 46940
rect 17568 46928 17574 46940
rect 17626 46928 17632 46980
rect 26584 46928 26590 46980
rect 26642 46928 26648 46980
rect 27136 46928 27142 46980
rect 27194 46968 27200 46980
rect 34039 46971 34097 46977
rect 34039 46968 34051 46971
rect 27194 46940 34051 46968
rect 27194 46928 27200 46940
rect 34039 46937 34051 46940
rect 34085 46937 34097 46971
rect 34039 46931 34097 46937
rect 1086 46810 58862 46832
rect 1086 46758 4228 46810
rect 4280 46758 4292 46810
rect 4344 46758 4356 46810
rect 4408 46758 4420 46810
rect 4472 46758 34948 46810
rect 35000 46758 35012 46810
rect 35064 46758 35076 46810
rect 35128 46758 35140 46810
rect 35192 46758 58862 46810
rect 1086 46736 58862 46758
rect 20512 46452 20518 46504
rect 20570 46492 20576 46504
rect 33763 46495 33821 46501
rect 33763 46492 33775 46495
rect 20570 46464 33775 46492
rect 20570 46452 20576 46464
rect 33763 46461 33775 46464
rect 33809 46461 33821 46495
rect 33763 46455 33821 46461
rect 55104 46452 55110 46504
rect 55162 46492 55168 46504
rect 58419 46495 58477 46501
rect 58419 46492 58431 46495
rect 55162 46464 58431 46492
rect 55162 46452 55168 46464
rect 58419 46461 58431 46464
rect 58465 46461 58477 46495
rect 58419 46455 58477 46461
rect 5424 46316 5430 46368
rect 5482 46356 5488 46368
rect 48023 46359 48081 46365
rect 48023 46356 48035 46359
rect 5482 46328 48035 46356
rect 5482 46316 5488 46328
rect 48023 46325 48035 46328
rect 48069 46325 48081 46359
rect 48023 46319 48081 46325
rect 1086 46266 58862 46288
rect 1086 46214 19588 46266
rect 19640 46214 19652 46266
rect 19704 46214 19716 46266
rect 19768 46214 19780 46266
rect 19832 46214 50308 46266
rect 50360 46214 50372 46266
rect 50424 46214 50436 46266
rect 50488 46214 50500 46266
rect 50552 46214 58862 46266
rect 1086 46192 58862 46214
rect 25940 46112 25946 46164
rect 25998 46152 26004 46164
rect 26124 46152 26130 46164
rect 25998 46124 26130 46152
rect 25998 46112 26004 46124
rect 26124 46112 26130 46124
rect 26182 46112 26188 46164
rect 2851 45883 2909 45889
rect 2851 45849 2863 45883
rect 2897 45880 2909 45883
rect 21340 45880 21346 45892
rect 2897 45852 21346 45880
rect 2897 45849 2909 45852
rect 2851 45843 2909 45849
rect 21340 45840 21346 45852
rect 21398 45840 21404 45892
rect 9196 45812 9202 45824
rect 9157 45784 9202 45812
rect 9196 45772 9202 45784
rect 9254 45772 9260 45824
rect 20512 45812 20518 45824
rect 20473 45784 20518 45812
rect 20512 45772 20518 45784
rect 20570 45772 20576 45824
rect 23180 45772 23186 45824
rect 23238 45812 23244 45824
rect 32935 45815 32993 45821
rect 32935 45812 32947 45815
rect 23238 45784 32947 45812
rect 23238 45772 23244 45784
rect 32935 45781 32947 45784
rect 32981 45781 32993 45815
rect 32935 45775 32993 45781
rect 1086 45722 58862 45744
rect 1086 45670 4228 45722
rect 4280 45670 4292 45722
rect 4344 45670 4356 45722
rect 4408 45670 4420 45722
rect 4472 45670 34948 45722
rect 35000 45670 35012 45722
rect 35064 45670 35076 45722
rect 35128 45670 35140 45722
rect 35192 45670 58862 45722
rect 1086 45648 58862 45670
rect 7448 45568 7454 45620
rect 7506 45608 7512 45620
rect 7724 45608 7730 45620
rect 7506 45580 7730 45608
rect 7506 45568 7512 45580
rect 7724 45568 7730 45580
rect 7782 45568 7788 45620
rect 7908 45568 7914 45620
rect 7966 45608 7972 45620
rect 20512 45608 20518 45620
rect 7966 45580 20518 45608
rect 7966 45568 7972 45580
rect 20512 45568 20518 45580
rect 20570 45568 20576 45620
rect 26216 45500 26222 45552
rect 26274 45540 26280 45552
rect 26584 45540 26590 45552
rect 26274 45512 26590 45540
rect 26274 45500 26280 45512
rect 26584 45500 26590 45512
rect 26642 45500 26648 45552
rect 38820 45500 38826 45552
rect 38878 45540 38884 45552
rect 39004 45540 39010 45552
rect 38878 45512 39010 45540
rect 38878 45500 38884 45512
rect 39004 45500 39010 45512
rect 39062 45500 39068 45552
rect 9564 45364 9570 45416
rect 9622 45404 9628 45416
rect 20975 45407 21033 45413
rect 20975 45404 20987 45407
rect 9622 45376 20987 45404
rect 9622 45364 9628 45376
rect 20975 45373 20987 45376
rect 21021 45373 21033 45407
rect 29436 45404 29442 45416
rect 29397 45376 29442 45404
rect 20975 45367 21033 45373
rect 29436 45364 29442 45376
rect 29494 45364 29500 45416
rect 39007 45407 39065 45413
rect 39007 45373 39019 45407
rect 39053 45373 39065 45407
rect 39007 45367 39065 45373
rect 17844 45296 17850 45348
rect 17902 45336 17908 45348
rect 39022 45336 39050 45367
rect 17902 45308 39050 45336
rect 17902 45296 17908 45308
rect 1086 45178 58862 45200
rect 1086 45126 19588 45178
rect 19640 45126 19652 45178
rect 19704 45126 19716 45178
rect 19768 45126 19780 45178
rect 19832 45126 50308 45178
rect 50360 45126 50372 45178
rect 50424 45126 50436 45178
rect 50488 45126 50500 45178
rect 50552 45126 58862 45178
rect 1086 45104 58862 45126
rect 16372 44684 16378 44736
rect 16430 44724 16436 44736
rect 36891 44727 36949 44733
rect 36891 44724 36903 44727
rect 16430 44696 36903 44724
rect 16430 44684 16436 44696
rect 36891 44693 36903 44696
rect 36937 44693 36949 44727
rect 36891 44687 36949 44693
rect 1086 44634 58862 44656
rect 1086 44582 4228 44634
rect 4280 44582 4292 44634
rect 4344 44582 4356 44634
rect 4408 44582 4420 44634
rect 4472 44582 34948 44634
rect 35000 44582 35012 44634
rect 35064 44582 35076 44634
rect 35128 44582 35140 44634
rect 35192 44582 58862 44634
rect 1086 44560 58862 44582
rect 13799 44387 13857 44393
rect 13799 44353 13811 44387
rect 13845 44384 13857 44387
rect 26860 44384 26866 44396
rect 13845 44356 26866 44384
rect 13845 44353 13857 44356
rect 13799 44347 13857 44353
rect 26860 44344 26866 44356
rect 26918 44344 26924 44396
rect 21910 44288 22122 44316
rect 5148 44208 5154 44260
rect 5206 44248 5212 44260
rect 21910 44248 21938 44288
rect 5206 44220 21938 44248
rect 22094 44248 22122 44288
rect 29896 44276 29902 44328
rect 29954 44316 29960 44328
rect 29991 44319 30049 44325
rect 29991 44316 30003 44319
rect 29954 44288 30003 44316
rect 29954 44276 29960 44288
rect 29991 44285 30003 44288
rect 30037 44285 30049 44319
rect 36612 44316 36618 44328
rect 36573 44288 36618 44316
rect 29991 44279 30049 44285
rect 36612 44276 36618 44288
rect 36670 44276 36676 44328
rect 38176 44316 38182 44328
rect 38137 44288 38182 44316
rect 38176 44276 38182 44288
rect 38234 44276 38240 44328
rect 42503 44319 42561 44325
rect 42503 44285 42515 44319
rect 42549 44285 42561 44319
rect 42503 44279 42561 44285
rect 42518 44248 42546 44279
rect 22094 44220 42546 44248
rect 5206 44208 5212 44220
rect 45536 44140 45542 44192
rect 45594 44180 45600 44192
rect 45720 44180 45726 44192
rect 45594 44152 45726 44180
rect 45594 44140 45600 44152
rect 45720 44140 45726 44152
rect 45778 44140 45784 44192
rect 1086 44090 58862 44112
rect 1086 44038 19588 44090
rect 19640 44038 19652 44090
rect 19704 44038 19716 44090
rect 19768 44038 19780 44090
rect 19832 44038 50308 44090
rect 50360 44038 50372 44090
rect 50424 44038 50436 44090
rect 50488 44038 50500 44090
rect 50552 44038 58862 44090
rect 1086 44016 58862 44038
rect 44892 43976 44898 43988
rect 44853 43948 44898 43976
rect 44892 43936 44898 43948
rect 44950 43936 44956 43988
rect 48296 43936 48302 43988
rect 48354 43976 48360 43988
rect 48354 43948 53126 43976
rect 48354 43936 48360 43948
rect 44803 43843 44861 43849
rect 44803 43809 44815 43843
rect 44849 43840 44861 43843
rect 48296 43840 48302 43852
rect 44849 43812 48302 43840
rect 44849 43809 44861 43812
rect 44803 43803 44861 43809
rect 48296 43800 48302 43812
rect 48354 43800 48360 43852
rect 52991 43843 53049 43849
rect 52991 43809 53003 43843
rect 53037 43840 53049 43843
rect 53098 43840 53126 43948
rect 53037 43812 53126 43840
rect 53037 43809 53049 43812
rect 52991 43803 53049 43809
rect 37440 43772 37446 43784
rect 37401 43744 37446 43772
rect 37440 43732 37446 43744
rect 37498 43732 37504 43784
rect 50964 43772 50970 43784
rect 48222 43744 50970 43772
rect 30264 43664 30270 43716
rect 30322 43704 30328 43716
rect 48222 43704 48250 43744
rect 50964 43732 50970 43744
rect 51022 43732 51028 43784
rect 51056 43732 51062 43784
rect 51114 43772 51120 43784
rect 51979 43775 52037 43781
rect 51979 43772 51991 43775
rect 51114 43744 51991 43772
rect 51114 43732 51120 43744
rect 51979 43741 51991 43744
rect 52025 43741 52037 43775
rect 51979 43735 52037 43741
rect 30322 43676 48250 43704
rect 30322 43664 30328 43676
rect 6715 43639 6773 43645
rect 6715 43605 6727 43639
rect 6761 43636 6773 43639
rect 20052 43636 20058 43648
rect 6761 43608 20058 43636
rect 6761 43605 6773 43608
rect 6715 43599 6773 43605
rect 20052 43596 20058 43608
rect 20110 43596 20116 43648
rect 23364 43596 23370 43648
rect 23422 43636 23428 43648
rect 44803 43639 44861 43645
rect 44803 43636 44815 43639
rect 23422 43608 44815 43636
rect 23422 43596 23428 43608
rect 44803 43605 44815 43608
rect 44849 43605 44861 43639
rect 44803 43599 44861 43605
rect 1086 43546 58862 43568
rect 1086 43494 4228 43546
rect 4280 43494 4292 43546
rect 4344 43494 4356 43546
rect 4408 43494 4420 43546
rect 4472 43494 34948 43546
rect 35000 43494 35012 43546
rect 35064 43494 35076 43546
rect 35128 43494 35140 43546
rect 35192 43494 58862 43546
rect 1086 43472 58862 43494
rect 14992 43432 14998 43444
rect 14953 43404 14998 43432
rect 14992 43392 14998 43404
rect 15050 43392 15056 43444
rect 34588 43324 34594 43376
rect 34646 43364 34652 43376
rect 34772 43364 34778 43376
rect 34646 43336 34778 43364
rect 34646 43324 34652 43336
rect 34772 43324 34778 43336
rect 34830 43324 34836 43376
rect 1379 43163 1437 43169
rect 1379 43129 1391 43163
rect 1425 43160 1437 43163
rect 20144 43160 20150 43172
rect 1425 43132 20150 43160
rect 1425 43129 1437 43132
rect 1379 43123 1437 43129
rect 20144 43120 20150 43132
rect 20202 43120 20208 43172
rect 9935 43095 9993 43101
rect 9935 43061 9947 43095
rect 9981 43092 9993 43095
rect 33852 43092 33858 43104
rect 9981 43064 33858 43092
rect 9981 43061 9993 43064
rect 9935 43055 9993 43061
rect 33852 43052 33858 43064
rect 33910 43052 33916 43104
rect 1086 43002 58862 43024
rect 1086 42950 19588 43002
rect 19640 42950 19652 43002
rect 19704 42950 19716 43002
rect 19768 42950 19780 43002
rect 19832 42950 50308 43002
rect 50360 42950 50372 43002
rect 50424 42950 50436 43002
rect 50488 42950 50500 43002
rect 50552 42950 58862 43002
rect 1086 42928 58862 42950
rect 1086 42458 58862 42480
rect 1086 42406 4228 42458
rect 4280 42406 4292 42458
rect 4344 42406 4356 42458
rect 4408 42406 4420 42458
rect 4472 42406 34948 42458
rect 35000 42406 35012 42458
rect 35064 42406 35076 42458
rect 35128 42406 35140 42458
rect 35192 42406 58862 42458
rect 1086 42384 58862 42406
rect 9932 42208 9938 42220
rect 9893 42180 9938 42208
rect 9932 42168 9938 42180
rect 9990 42168 9996 42220
rect 13520 42100 13526 42152
rect 13578 42140 13584 42152
rect 36063 42143 36121 42149
rect 36063 42140 36075 42143
rect 13578 42112 36075 42140
rect 13578 42100 13584 42112
rect 36063 42109 36075 42112
rect 36109 42109 36121 42143
rect 36063 42103 36121 42109
rect 1086 41914 58862 41936
rect 1086 41862 19588 41914
rect 19640 41862 19652 41914
rect 19704 41862 19716 41914
rect 19768 41862 19780 41914
rect 19832 41862 50308 41914
rect 50360 41862 50372 41914
rect 50424 41862 50436 41914
rect 50488 41862 50500 41914
rect 50552 41862 58862 41914
rect 1086 41840 58862 41862
rect 1086 41370 58862 41392
rect 1086 41318 4228 41370
rect 4280 41318 4292 41370
rect 4344 41318 4356 41370
rect 4408 41318 4420 41370
rect 4472 41318 34948 41370
rect 35000 41318 35012 41370
rect 35064 41318 35076 41370
rect 35128 41318 35140 41370
rect 35192 41318 58862 41370
rect 1086 41296 58862 41318
rect 19960 41256 19966 41268
rect 19921 41228 19966 41256
rect 19960 41216 19966 41228
rect 20018 41216 20024 41268
rect 7543 41055 7601 41061
rect 7543 41021 7555 41055
rect 7589 41021 7601 41055
rect 7543 41015 7601 41021
rect 11131 41055 11189 41061
rect 11131 41021 11143 41055
rect 11177 41052 11189 41055
rect 28332 41052 28338 41064
rect 11177 41024 28338 41052
rect 11177 41021 11189 41024
rect 11131 41015 11189 41021
rect 7558 40984 7586 41015
rect 28332 41012 28338 41024
rect 28390 41012 28396 41064
rect 24192 40984 24198 40996
rect 7558 40956 24198 40984
rect 24192 40944 24198 40956
rect 24250 40944 24256 40996
rect 1086 40826 58862 40848
rect 1086 40774 19588 40826
rect 19640 40774 19652 40826
rect 19704 40774 19716 40826
rect 19768 40774 19780 40826
rect 19832 40774 50308 40826
rect 50360 40774 50372 40826
rect 50424 40774 50436 40826
rect 50488 40774 50500 40826
rect 50552 40774 58862 40826
rect 1086 40752 58862 40774
rect 6439 40375 6497 40381
rect 6439 40341 6451 40375
rect 6485 40372 6497 40375
rect 27136 40372 27142 40384
rect 6485 40344 27142 40372
rect 6485 40341 6497 40344
rect 6439 40335 6497 40341
rect 27136 40332 27142 40344
rect 27194 40332 27200 40384
rect 50964 40332 50970 40384
rect 51022 40372 51028 40384
rect 55935 40375 55993 40381
rect 55935 40372 55947 40375
rect 51022 40344 55947 40372
rect 51022 40332 51028 40344
rect 55935 40341 55947 40344
rect 55981 40341 55993 40375
rect 55935 40335 55993 40341
rect 1086 40282 58862 40304
rect 1086 40230 4228 40282
rect 4280 40230 4292 40282
rect 4344 40230 4356 40282
rect 4408 40230 4420 40282
rect 4472 40230 34948 40282
rect 35000 40230 35012 40282
rect 35064 40230 35076 40282
rect 35128 40230 35140 40282
rect 35192 40230 58862 40282
rect 1086 40208 58862 40230
rect 4964 40100 4970 40112
rect 4925 40072 4970 40100
rect 4964 40060 4970 40072
rect 5022 40060 5028 40112
rect 14624 40100 14630 40112
rect 14585 40072 14630 40100
rect 14624 40060 14630 40072
rect 14682 40060 14688 40112
rect 28792 40060 28798 40112
rect 28850 40100 28856 40112
rect 57591 40103 57649 40109
rect 57591 40100 57603 40103
rect 28850 40072 57603 40100
rect 28850 40060 28856 40072
rect 57591 40069 57603 40072
rect 57637 40069 57649 40103
rect 57591 40063 57649 40069
rect 1086 39738 58862 39760
rect 1086 39686 19588 39738
rect 19640 39686 19652 39738
rect 19704 39686 19716 39738
rect 19768 39686 19780 39738
rect 19832 39686 50308 39738
rect 50360 39686 50372 39738
rect 50424 39686 50436 39738
rect 50488 39686 50500 39738
rect 50552 39686 58862 39738
rect 1086 39664 58862 39686
rect 20512 39380 20518 39432
rect 20570 39420 20576 39432
rect 23364 39420 23370 39432
rect 20570 39392 23370 39420
rect 20570 39380 20576 39392
rect 23364 39380 23370 39392
rect 23422 39380 23428 39432
rect 27504 39380 27510 39432
rect 27562 39420 27568 39432
rect 41859 39423 41917 39429
rect 41859 39420 41871 39423
rect 27562 39392 41871 39420
rect 27562 39380 27568 39392
rect 41859 39389 41871 39392
rect 41905 39389 41917 39423
rect 41859 39383 41917 39389
rect 7356 39312 7362 39364
rect 7414 39352 7420 39364
rect 7540 39352 7546 39364
rect 7414 39324 7546 39352
rect 7414 39312 7420 39324
rect 7540 39312 7546 39324
rect 7598 39312 7604 39364
rect 5240 39244 5246 39296
rect 5298 39284 5304 39296
rect 21803 39287 21861 39293
rect 21803 39284 21815 39287
rect 5298 39256 21815 39284
rect 5298 39244 5304 39256
rect 21803 39253 21815 39256
rect 21849 39253 21861 39287
rect 36980 39284 36986 39296
rect 36941 39256 36986 39284
rect 21803 39247 21861 39253
rect 36980 39244 36986 39256
rect 37038 39244 37044 39296
rect 49584 39244 49590 39296
rect 49642 39284 49648 39296
rect 56119 39287 56177 39293
rect 56119 39284 56131 39287
rect 49642 39256 56131 39284
rect 49642 39244 49648 39256
rect 56119 39253 56131 39256
rect 56165 39253 56177 39287
rect 56119 39247 56177 39253
rect 1086 39194 58862 39216
rect 1086 39142 4228 39194
rect 4280 39142 4292 39194
rect 4344 39142 4356 39194
rect 4408 39142 4420 39194
rect 4472 39142 34948 39194
rect 35000 39142 35012 39194
rect 35064 39142 35076 39194
rect 35128 39142 35140 39194
rect 35192 39142 58862 39194
rect 1086 39120 58862 39142
rect 19132 39040 19138 39092
rect 19190 39080 19196 39092
rect 23183 39083 23241 39089
rect 23183 39080 23195 39083
rect 19190 39052 23195 39080
rect 19190 39040 19196 39052
rect 23183 39049 23195 39052
rect 23229 39049 23241 39083
rect 23183 39043 23241 39049
rect 1086 38650 58862 38672
rect 1086 38598 19588 38650
rect 19640 38598 19652 38650
rect 19704 38598 19716 38650
rect 19768 38598 19780 38650
rect 19832 38598 50308 38650
rect 50360 38598 50372 38650
rect 50424 38598 50436 38650
rect 50488 38598 50500 38650
rect 50552 38598 58862 38650
rect 1086 38576 58862 38598
rect 26679 38199 26737 38205
rect 26679 38165 26691 38199
rect 26725 38196 26737 38199
rect 28976 38196 28982 38208
rect 26725 38168 28982 38196
rect 26725 38165 26737 38168
rect 26679 38159 26737 38165
rect 28976 38156 28982 38168
rect 29034 38156 29040 38208
rect 1086 38106 58862 38128
rect 1086 38054 4228 38106
rect 4280 38054 4292 38106
rect 4344 38054 4356 38106
rect 4408 38054 4420 38106
rect 4472 38054 34948 38106
rect 35000 38054 35012 38106
rect 35064 38054 35076 38106
rect 35128 38054 35140 38106
rect 35192 38054 58862 38106
rect 1086 38032 58862 38054
rect 1086 37562 58862 37584
rect 1086 37510 19588 37562
rect 19640 37510 19652 37562
rect 19704 37510 19716 37562
rect 19768 37510 19780 37562
rect 19832 37510 50308 37562
rect 50360 37510 50372 37562
rect 50424 37510 50436 37562
rect 50488 37510 50500 37562
rect 50552 37510 58862 37562
rect 1086 37488 58862 37510
rect 21800 37448 21806 37460
rect 21761 37420 21806 37448
rect 21800 37408 21806 37420
rect 21858 37408 21864 37460
rect 8644 37272 8650 37324
rect 8702 37312 8708 37324
rect 8736 37312 8742 37324
rect 8702 37284 8742 37312
rect 8702 37272 8708 37284
rect 8736 37272 8742 37284
rect 8794 37272 8800 37324
rect 29896 37272 29902 37324
rect 29954 37312 29960 37324
rect 29988 37312 29994 37324
rect 29954 37284 29994 37312
rect 29954 37272 29960 37284
rect 29988 37272 29994 37284
rect 30046 37272 30052 37324
rect 37440 37272 37446 37324
rect 37498 37312 37504 37324
rect 46272 37312 46278 37324
rect 37498 37284 46278 37312
rect 37498 37272 37504 37284
rect 46272 37272 46278 37284
rect 46330 37272 46336 37324
rect 6804 37204 6810 37256
rect 6862 37244 6868 37256
rect 6862 37216 11358 37244
rect 6862 37204 6868 37216
rect 11330 37176 11358 37216
rect 25299 37179 25357 37185
rect 25299 37176 25311 37179
rect 4706 37148 11266 37176
rect 11330 37148 25311 37176
rect 1100 37068 1106 37120
rect 1158 37108 1164 37120
rect 4706 37108 4734 37148
rect 11128 37108 11134 37120
rect 1158 37080 4734 37108
rect 11089 37080 11134 37108
rect 1158 37068 1164 37080
rect 11128 37068 11134 37080
rect 11186 37068 11192 37120
rect 11238 37108 11266 37148
rect 25299 37145 25311 37148
rect 25345 37145 25357 37179
rect 25299 37139 25357 37145
rect 26955 37111 27013 37117
rect 26955 37108 26967 37111
rect 11238 37080 26967 37108
rect 26955 37077 26967 37080
rect 27001 37077 27013 37111
rect 26955 37071 27013 37077
rect 38544 37068 38550 37120
rect 38602 37108 38608 37120
rect 45079 37111 45137 37117
rect 45079 37108 45091 37111
rect 38602 37080 45091 37108
rect 38602 37068 38608 37080
rect 45079 37077 45091 37080
rect 45125 37077 45137 37111
rect 45079 37071 45137 37077
rect 1086 37018 58862 37040
rect 1086 36966 4228 37018
rect 4280 36966 4292 37018
rect 4344 36966 4356 37018
rect 4408 36966 4420 37018
rect 4472 36966 34948 37018
rect 35000 36966 35012 37018
rect 35064 36966 35076 37018
rect 35128 36966 35140 37018
rect 35192 36966 58862 37018
rect 1086 36944 58862 36966
rect 19408 36904 19414 36916
rect 19369 36876 19414 36904
rect 19408 36864 19414 36876
rect 19466 36864 19472 36916
rect 34312 36728 34318 36780
rect 34370 36768 34376 36780
rect 53083 36771 53141 36777
rect 53083 36768 53095 36771
rect 34370 36740 53095 36768
rect 34370 36728 34376 36740
rect 53083 36737 53095 36740
rect 53129 36737 53141 36771
rect 53083 36731 53141 36737
rect 3768 36660 3774 36712
rect 3826 36700 3832 36712
rect 4691 36703 4749 36709
rect 4691 36700 4703 36703
rect 3826 36672 4703 36700
rect 3826 36660 3832 36672
rect 4691 36669 4703 36672
rect 4737 36669 4749 36703
rect 11772 36700 11778 36712
rect 11733 36672 11778 36700
rect 4691 36663 4749 36669
rect 11772 36660 11778 36672
rect 11830 36660 11836 36712
rect 15455 36703 15513 36709
rect 15455 36669 15467 36703
rect 15501 36669 15513 36703
rect 15455 36663 15513 36669
rect 35051 36703 35109 36709
rect 35051 36669 35063 36703
rect 35097 36700 35109 36703
rect 35232 36700 35238 36712
rect 35097 36672 35238 36700
rect 35097 36669 35109 36672
rect 35051 36663 35109 36669
rect 15470 36632 15498 36663
rect 35232 36660 35238 36672
rect 35290 36660 35296 36712
rect 40752 36632 40758 36644
rect 15470 36604 40758 36632
rect 40752 36592 40758 36604
rect 40810 36592 40816 36644
rect 1086 36474 58862 36496
rect 1086 36422 19588 36474
rect 19640 36422 19652 36474
rect 19704 36422 19716 36474
rect 19768 36422 19780 36474
rect 19832 36422 50308 36474
rect 50360 36422 50372 36474
rect 50424 36422 50436 36474
rect 50488 36422 50500 36474
rect 50552 36422 58862 36474
rect 1086 36400 58862 36422
rect 25940 36320 25946 36372
rect 25998 36360 26004 36372
rect 26124 36360 26130 36372
rect 25998 36332 26130 36360
rect 25998 36320 26004 36332
rect 26124 36320 26130 36332
rect 26182 36320 26188 36372
rect 6344 36020 6350 36032
rect 6305 35992 6350 36020
rect 6344 35980 6350 35992
rect 6402 35980 6408 36032
rect 26216 35980 26222 36032
rect 26274 36020 26280 36032
rect 26400 36020 26406 36032
rect 26274 35992 26406 36020
rect 26274 35980 26280 35992
rect 26400 35980 26406 35992
rect 26458 35980 26464 36032
rect 38084 36020 38090 36032
rect 38045 35992 38090 36020
rect 38084 35980 38090 35992
rect 38142 35980 38148 36032
rect 1086 35930 58862 35952
rect 1086 35878 4228 35930
rect 4280 35878 4292 35930
rect 4344 35878 4356 35930
rect 4408 35878 4420 35930
rect 4472 35878 34948 35930
rect 35000 35878 35012 35930
rect 35064 35878 35076 35930
rect 35128 35878 35140 35930
rect 35192 35878 58862 35930
rect 1086 35856 58862 35878
rect 38360 35816 38366 35828
rect 38321 35788 38366 35816
rect 38360 35776 38366 35788
rect 38418 35776 38424 35828
rect 4507 35615 4565 35621
rect 4507 35581 4519 35615
rect 4553 35612 4565 35615
rect 21432 35612 21438 35624
rect 4553 35584 21438 35612
rect 4553 35581 4565 35584
rect 4507 35575 4565 35581
rect 21432 35572 21438 35584
rect 21490 35572 21496 35624
rect 55656 35612 55662 35624
rect 55617 35584 55662 35612
rect 55656 35572 55662 35584
rect 55714 35572 55720 35624
rect 1086 35386 58862 35408
rect 1086 35334 19588 35386
rect 19640 35334 19652 35386
rect 19704 35334 19716 35386
rect 19768 35334 19780 35386
rect 19832 35334 50308 35386
rect 50360 35334 50372 35386
rect 50424 35334 50436 35386
rect 50488 35334 50500 35386
rect 50552 35334 58862 35386
rect 1086 35312 58862 35334
rect 1100 34892 1106 34944
rect 1158 34932 1164 34944
rect 16283 34935 16341 34941
rect 16283 34932 16295 34935
rect 1158 34904 16295 34932
rect 1158 34892 1164 34904
rect 16283 34901 16295 34904
rect 16329 34901 16341 34935
rect 16283 34895 16341 34901
rect 1086 34842 58862 34864
rect 1086 34790 4228 34842
rect 4280 34790 4292 34842
rect 4344 34790 4356 34842
rect 4408 34790 4420 34842
rect 4472 34790 34948 34842
rect 35000 34790 35012 34842
rect 35064 34790 35076 34842
rect 35128 34790 35140 34842
rect 35192 34790 58862 34842
rect 1086 34768 58862 34790
rect 7356 34484 7362 34536
rect 7414 34524 7420 34536
rect 7632 34524 7638 34536
rect 7414 34496 7638 34524
rect 7414 34484 7420 34496
rect 7632 34484 7638 34496
rect 7690 34484 7696 34536
rect 22996 34484 23002 34536
rect 23054 34524 23060 34536
rect 23180 34524 23186 34536
rect 23054 34496 23186 34524
rect 23054 34484 23060 34496
rect 23180 34484 23186 34496
rect 23238 34484 23244 34536
rect 43055 34527 43113 34533
rect 43055 34493 43067 34527
rect 43101 34524 43113 34527
rect 44984 34524 44990 34536
rect 43101 34496 44990 34524
rect 43101 34493 43113 34496
rect 43055 34487 43113 34493
rect 44984 34484 44990 34496
rect 45042 34484 45048 34536
rect 1086 34298 58862 34320
rect 1086 34246 19588 34298
rect 19640 34246 19652 34298
rect 19704 34246 19716 34298
rect 19768 34246 19780 34298
rect 19832 34246 50308 34298
rect 50360 34246 50372 34298
rect 50424 34246 50436 34298
rect 50488 34246 50500 34298
rect 50552 34246 58862 34298
rect 1086 34224 58862 34246
rect 6623 33847 6681 33853
rect 6623 33813 6635 33847
rect 6669 33844 6681 33847
rect 42040 33844 42046 33856
rect 6669 33816 42046 33844
rect 6669 33813 6681 33816
rect 6623 33807 6681 33813
rect 42040 33804 42046 33816
rect 42098 33804 42104 33856
rect 48480 33804 48486 33856
rect 48538 33844 48544 33856
rect 48664 33844 48670 33856
rect 48538 33816 48670 33844
rect 48538 33804 48544 33816
rect 48664 33804 48670 33816
rect 48722 33804 48728 33856
rect 1086 33754 58862 33776
rect 1086 33702 4228 33754
rect 4280 33702 4292 33754
rect 4344 33702 4356 33754
rect 4408 33702 4420 33754
rect 4472 33702 34948 33754
rect 35000 33702 35012 33754
rect 35064 33702 35076 33754
rect 35128 33702 35140 33754
rect 35192 33702 58862 33754
rect 1086 33680 58862 33702
rect 1086 33210 58862 33232
rect 1086 33158 19588 33210
rect 19640 33158 19652 33210
rect 19704 33158 19716 33210
rect 19768 33158 19780 33210
rect 19832 33158 50308 33210
rect 50360 33158 50372 33210
rect 50424 33158 50436 33210
rect 50488 33158 50500 33210
rect 50552 33158 58862 33210
rect 1086 33136 58862 33158
rect 22628 32960 22634 32972
rect 19150 32932 22634 32960
rect 4323 32895 4381 32901
rect 4323 32861 4335 32895
rect 4369 32892 4381 32895
rect 19150 32892 19178 32932
rect 22628 32920 22634 32932
rect 22686 32920 22692 32972
rect 4369 32864 19178 32892
rect 4369 32861 4381 32864
rect 4323 32855 4381 32861
rect 9196 32716 9202 32768
rect 9254 32756 9260 32768
rect 9472 32756 9478 32768
rect 9254 32728 9478 32756
rect 9254 32716 9260 32728
rect 9472 32716 9478 32728
rect 9530 32716 9536 32768
rect 11864 32756 11870 32768
rect 11825 32728 11870 32756
rect 11864 32716 11870 32728
rect 11922 32716 11928 32768
rect 22628 32716 22634 32768
rect 22686 32756 22692 32768
rect 32472 32756 32478 32768
rect 22686 32728 32478 32756
rect 22686 32716 22692 32728
rect 32472 32716 32478 32728
rect 32530 32716 32536 32768
rect 1086 32666 58862 32688
rect 1086 32614 4228 32666
rect 4280 32614 4292 32666
rect 4344 32614 4356 32666
rect 4408 32614 4420 32666
rect 4472 32614 34948 32666
rect 35000 32614 35012 32666
rect 35064 32614 35076 32666
rect 35128 32614 35140 32666
rect 35192 32614 58862 32666
rect 1086 32592 58862 32614
rect 2480 32512 2486 32564
rect 2538 32552 2544 32564
rect 11864 32552 11870 32564
rect 2538 32524 11870 32552
rect 2538 32512 2544 32524
rect 11864 32512 11870 32524
rect 11922 32512 11928 32564
rect 23180 32444 23186 32496
rect 23238 32484 23244 32496
rect 23548 32484 23554 32496
rect 23238 32456 23554 32484
rect 23238 32444 23244 32456
rect 23548 32444 23554 32456
rect 23606 32444 23612 32496
rect 8736 32376 8742 32428
rect 8794 32416 8800 32428
rect 9196 32416 9202 32428
rect 8794 32388 9202 32416
rect 8794 32376 8800 32388
rect 9196 32376 9202 32388
rect 9254 32376 9260 32428
rect 26952 32376 26958 32428
rect 27010 32416 27016 32428
rect 27136 32416 27142 32428
rect 27010 32388 27142 32416
rect 27010 32376 27016 32388
rect 27136 32376 27142 32388
rect 27194 32376 27200 32428
rect 1086 32122 58862 32144
rect 1086 32070 19588 32122
rect 19640 32070 19652 32122
rect 19704 32070 19716 32122
rect 19768 32070 19780 32122
rect 19832 32070 50308 32122
rect 50360 32070 50372 32122
rect 50424 32070 50436 32122
rect 50488 32070 50500 32122
rect 50552 32070 58862 32122
rect 1086 32048 58862 32070
rect 21984 31764 21990 31816
rect 22042 31804 22048 31816
rect 54739 31807 54797 31813
rect 54739 31804 54751 31807
rect 22042 31776 54751 31804
rect 22042 31764 22048 31776
rect 54739 31773 54751 31776
rect 54785 31773 54797 31807
rect 54739 31767 54797 31773
rect 1086 31578 58862 31600
rect 1086 31526 4228 31578
rect 4280 31526 4292 31578
rect 4344 31526 4356 31578
rect 4408 31526 4420 31578
rect 4472 31526 34948 31578
rect 35000 31526 35012 31578
rect 35064 31526 35076 31578
rect 35128 31526 35140 31578
rect 35192 31526 58862 31578
rect 1086 31504 58862 31526
rect 8736 31260 8742 31272
rect 8616 31232 8742 31260
rect 8616 31178 8644 31232
rect 8736 31220 8742 31232
rect 8794 31220 8800 31272
rect 11036 31260 11042 31272
rect 9182 31232 11042 31260
rect 11036 31220 11042 31232
rect 11094 31220 11100 31272
rect 11220 31260 11226 31272
rect 11181 31232 11226 31260
rect 11220 31220 11226 31232
rect 11278 31220 11284 31272
rect 36063 31263 36121 31269
rect 36063 31229 36075 31263
rect 36109 31260 36121 31263
rect 38820 31260 38826 31272
rect 36109 31232 38826 31260
rect 36109 31229 36121 31232
rect 36063 31223 36121 31229
rect 38820 31220 38826 31232
rect 38878 31220 38884 31272
rect 8828 31084 8834 31136
rect 8886 31084 8892 31136
rect 9012 31084 9018 31136
rect 9070 31124 9076 31136
rect 28424 31124 28430 31136
rect 9070 31096 28430 31124
rect 9070 31084 9076 31096
rect 28424 31084 28430 31096
rect 28482 31084 28488 31136
rect 1086 31034 58862 31056
rect 1086 30982 19588 31034
rect 19640 30982 19652 31034
rect 19704 30982 19716 31034
rect 19768 30982 19780 31034
rect 19832 30982 50308 31034
rect 50360 30982 50372 31034
rect 50424 30982 50436 31034
rect 50488 30982 50500 31034
rect 50552 30982 58862 31034
rect 1086 30960 58862 30982
rect 11036 30880 11042 30932
rect 11094 30920 11100 30932
rect 27872 30920 27878 30932
rect 11094 30892 27878 30920
rect 11094 30880 11100 30892
rect 27872 30880 27878 30892
rect 27930 30880 27936 30932
rect 8736 30812 8742 30864
rect 8794 30852 8800 30864
rect 28700 30852 28706 30864
rect 8794 30824 28706 30852
rect 8794 30812 8800 30824
rect 28700 30812 28706 30824
rect 28758 30812 28764 30864
rect 1086 30490 58862 30512
rect 1086 30438 4228 30490
rect 4280 30438 4292 30490
rect 4344 30438 4356 30490
rect 4408 30438 4420 30490
rect 4472 30438 34948 30490
rect 35000 30438 35012 30490
rect 35064 30438 35076 30490
rect 35128 30438 35140 30490
rect 35192 30438 58862 30490
rect 1086 30416 58862 30438
rect 54003 30243 54061 30249
rect 54003 30209 54015 30243
rect 54049 30240 54061 30243
rect 54049 30212 54138 30240
rect 54049 30209 54061 30212
rect 54003 30203 54061 30209
rect 8460 30132 8466 30184
rect 8518 30132 8524 30184
rect 13152 30172 13158 30184
rect 9182 30144 13158 30172
rect 13152 30132 13158 30144
rect 13210 30132 13216 30184
rect 14992 30132 14998 30184
rect 15050 30172 15056 30184
rect 17111 30175 17169 30181
rect 17111 30172 17123 30175
rect 15050 30144 17123 30172
rect 15050 30132 15056 30144
rect 17111 30141 17123 30144
rect 17157 30141 17169 30175
rect 17111 30135 17169 30141
rect 29439 30175 29497 30181
rect 29439 30141 29451 30175
rect 29485 30172 29497 30175
rect 29528 30172 29534 30184
rect 29485 30144 29534 30172
rect 29485 30141 29497 30144
rect 29439 30135 29497 30141
rect 29528 30132 29534 30144
rect 29586 30132 29592 30184
rect 48112 30172 48118 30184
rect 48073 30144 48118 30172
rect 48112 30132 48118 30144
rect 48170 30132 48176 30184
rect 48480 30172 48486 30184
rect 48441 30144 48486 30172
rect 48480 30132 48486 30144
rect 48538 30132 48544 30184
rect 8478 30056 8506 30132
rect 39924 30064 39930 30116
rect 39982 30104 39988 30116
rect 54110 30104 54138 30212
rect 39982 30076 54138 30104
rect 39982 30064 39988 30076
rect 8828 29996 8834 30048
rect 8886 29996 8892 30048
rect 9012 29996 9018 30048
rect 9070 30036 9076 30048
rect 25480 30036 25486 30048
rect 9070 30008 25486 30036
rect 9070 29996 9076 30008
rect 25480 29996 25486 30008
rect 25538 29996 25544 30048
rect 1086 29946 58862 29968
rect 1086 29894 19588 29946
rect 19640 29894 19652 29946
rect 19704 29894 19716 29946
rect 19768 29894 19780 29946
rect 19832 29894 50308 29946
rect 50360 29894 50372 29946
rect 50424 29894 50436 29946
rect 50488 29894 50500 29946
rect 50552 29894 58862 29946
rect 1086 29872 58862 29894
rect 13152 29792 13158 29844
rect 13210 29832 13216 29844
rect 27228 29832 27234 29844
rect 13210 29804 27234 29832
rect 13210 29792 13216 29804
rect 27228 29792 27234 29804
rect 27286 29792 27292 29844
rect 1008 29724 1014 29776
rect 1066 29764 1072 29776
rect 48480 29764 48486 29776
rect 1066 29736 48486 29764
rect 1066 29724 1072 29736
rect 48480 29724 48486 29736
rect 48538 29724 48544 29776
rect 7724 29656 7730 29708
rect 7782 29696 7788 29708
rect 48112 29696 48118 29708
rect 7782 29668 48118 29696
rect 7782 29656 7788 29668
rect 48112 29656 48118 29668
rect 48170 29656 48176 29708
rect 8460 29588 8466 29640
rect 8518 29628 8524 29640
rect 27688 29628 27694 29640
rect 8518 29600 27694 29628
rect 8518 29588 8524 29600
rect 27688 29588 27694 29600
rect 27746 29588 27752 29640
rect 8828 29520 8834 29572
rect 8886 29560 8892 29572
rect 25848 29560 25854 29572
rect 8886 29532 25854 29560
rect 8886 29520 8892 29532
rect 25848 29520 25854 29532
rect 25906 29520 25912 29572
rect 15636 29492 15642 29504
rect 15597 29464 15642 29492
rect 15636 29452 15642 29464
rect 15694 29452 15700 29504
rect 1086 29402 58862 29424
rect 1086 29350 4228 29402
rect 4280 29350 4292 29402
rect 4344 29350 4356 29402
rect 4408 29350 4420 29402
rect 4472 29350 34948 29402
rect 35000 29350 35012 29402
rect 35064 29350 35076 29402
rect 35128 29350 35140 29402
rect 35192 29350 58862 29402
rect 1086 29328 58862 29350
rect 3587 29291 3645 29297
rect 3587 29257 3599 29291
rect 3633 29288 3645 29291
rect 27136 29288 27142 29300
rect 3633 29260 27142 29288
rect 3633 29257 3645 29260
rect 3587 29251 3645 29257
rect 27136 29248 27142 29260
rect 27194 29248 27200 29300
rect 8828 29152 8834 29164
rect 8800 29112 8834 29152
rect 8886 29112 8892 29164
rect 26308 29152 26314 29164
rect 8998 29124 26314 29152
rect 26308 29112 26314 29124
rect 26366 29112 26372 29164
rect 8800 29070 8828 29112
rect 12048 29044 12054 29096
rect 12106 29084 12112 29096
rect 30359 29087 30417 29093
rect 30359 29084 30371 29087
rect 12106 29056 30371 29084
rect 12106 29044 12112 29056
rect 30359 29053 30371 29056
rect 30405 29053 30417 29087
rect 30359 29047 30417 29053
rect 19040 28976 19046 29028
rect 19098 29016 19104 29028
rect 19132 29016 19138 29028
rect 19098 28988 19138 29016
rect 19098 28976 19104 28988
rect 19132 28976 19138 28988
rect 19190 28976 19196 29028
rect 24008 28976 24014 29028
rect 24066 29016 24072 29028
rect 24100 29016 24106 29028
rect 24066 28988 24106 29016
rect 24066 28976 24072 28988
rect 24100 28976 24106 28988
rect 24158 28976 24164 29028
rect 34680 28976 34686 29028
rect 34738 29016 34744 29028
rect 34772 29016 34778 29028
rect 34738 28988 34778 29016
rect 34738 28976 34744 28988
rect 34772 28976 34778 28988
rect 34830 28976 34836 29028
rect 48296 28976 48302 29028
rect 48354 29016 48360 29028
rect 48664 29016 48670 29028
rect 48354 28988 48670 29016
rect 48354 28976 48360 28988
rect 48664 28976 48670 28988
rect 48722 28976 48728 29028
rect 24376 28948 24382 28960
rect 8722 28920 24382 28948
rect 24376 28908 24382 28920
rect 24434 28908 24440 28960
rect 1086 28858 58862 28880
rect 1086 28806 19588 28858
rect 19640 28806 19652 28858
rect 19704 28806 19716 28858
rect 19768 28806 19780 28858
rect 19832 28806 50308 28858
rect 50360 28806 50372 28858
rect 50424 28806 50436 28858
rect 50488 28806 50500 28858
rect 50552 28806 58862 28858
rect 1086 28784 58862 28806
rect 27596 28744 27602 28756
rect 27557 28716 27602 28744
rect 27596 28704 27602 28716
rect 27654 28704 27660 28756
rect 23272 28636 23278 28688
rect 23330 28676 23336 28688
rect 23456 28676 23462 28688
rect 23330 28648 23462 28676
rect 23330 28636 23336 28648
rect 23456 28636 23462 28648
rect 23514 28636 23520 28688
rect 3676 28364 3682 28416
rect 3734 28404 3740 28416
rect 25943 28407 26001 28413
rect 25943 28404 25955 28407
rect 3734 28376 25955 28404
rect 3734 28364 3740 28376
rect 25943 28373 25955 28376
rect 25989 28373 26001 28407
rect 34772 28404 34778 28416
rect 34733 28376 34778 28404
rect 25943 28367 26001 28373
rect 34772 28364 34778 28376
rect 34830 28364 34836 28416
rect 1086 28314 58862 28336
rect 1086 28262 4228 28314
rect 4280 28262 4292 28314
rect 4344 28262 4356 28314
rect 4408 28262 4420 28314
rect 4472 28262 34948 28314
rect 35000 28262 35012 28314
rect 35064 28262 35076 28314
rect 35128 28262 35140 28314
rect 35192 28262 58862 28314
rect 1086 28240 58862 28262
rect 13888 28160 13894 28212
rect 13946 28200 13952 28212
rect 34772 28200 34778 28212
rect 13946 28172 34778 28200
rect 13946 28160 13952 28172
rect 34772 28160 34778 28172
rect 34830 28160 34836 28212
rect 8552 28064 8558 28076
rect 8446 28036 8558 28064
rect 8552 28024 8558 28036
rect 8610 28024 8616 28076
rect 8920 28024 8926 28076
rect 8978 28064 8984 28076
rect 25388 28064 25394 28076
rect 8978 28036 25394 28064
rect 8978 28024 8984 28036
rect 25388 28024 25394 28036
rect 25446 28024 25452 28076
rect 8828 27956 8834 28008
rect 8886 27996 8892 28008
rect 24284 27996 24290 28008
rect 8886 27968 24290 27996
rect 8886 27956 8892 27968
rect 24284 27956 24290 27968
rect 24342 27956 24348 28008
rect 37808 27996 37814 28008
rect 37769 27968 37814 27996
rect 37808 27956 37814 27968
rect 37866 27956 37872 28008
rect 8478 27860 8506 27948
rect 8552 27860 8558 27872
rect 8478 27832 8558 27860
rect 8552 27820 8558 27832
rect 8610 27820 8616 27872
rect 22812 27860 22818 27872
rect 8722 27832 22818 27860
rect 22812 27820 22818 27832
rect 22870 27820 22876 27872
rect 1086 27770 58862 27792
rect 1086 27718 19588 27770
rect 19640 27718 19652 27770
rect 19704 27718 19716 27770
rect 19768 27718 19780 27770
rect 19832 27718 50308 27770
rect 50360 27718 50372 27770
rect 50424 27718 50436 27770
rect 50488 27718 50500 27770
rect 50552 27718 58862 27770
rect 1086 27696 58862 27718
rect 9288 27616 9294 27668
rect 9346 27656 9352 27668
rect 9472 27656 9478 27668
rect 9346 27628 9478 27656
rect 9346 27616 9352 27628
rect 9472 27616 9478 27628
rect 9530 27616 9536 27668
rect 13336 27616 13342 27668
rect 13394 27656 13400 27668
rect 13888 27656 13894 27668
rect 13394 27628 13894 27656
rect 13394 27616 13400 27628
rect 13888 27616 13894 27628
rect 13946 27616 13952 27668
rect 26400 27616 26406 27668
rect 26458 27656 26464 27668
rect 26492 27656 26498 27668
rect 26458 27628 26498 27656
rect 26458 27616 26464 27628
rect 26492 27616 26498 27628
rect 26550 27616 26556 27668
rect 28424 27616 28430 27668
rect 28482 27656 28488 27668
rect 29160 27656 29166 27668
rect 28482 27628 29166 27656
rect 28482 27616 28488 27628
rect 29160 27616 29166 27628
rect 29218 27616 29224 27668
rect 18856 27548 18862 27600
rect 18914 27588 18920 27600
rect 18948 27588 18954 27600
rect 18914 27560 18954 27588
rect 18914 27548 18920 27560
rect 18948 27548 18954 27560
rect 19006 27548 19012 27600
rect 1086 27226 58862 27248
rect 1086 27174 4228 27226
rect 4280 27174 4292 27226
rect 4344 27174 4356 27226
rect 4408 27174 4420 27226
rect 4472 27174 34948 27226
rect 35000 27174 35012 27226
rect 35064 27174 35076 27226
rect 35128 27174 35140 27226
rect 35192 27174 58862 27226
rect 1086 27152 58862 27174
rect 8414 26970 8420 27022
rect 8472 26970 8478 27022
rect 8828 27004 8834 27056
rect 8886 27044 8892 27056
rect 16556 27044 16562 27056
rect 8886 27016 16562 27044
rect 8886 27004 8892 27016
rect 16556 27004 16562 27016
rect 16614 27004 16620 27056
rect 8552 26908 8558 26920
rect 8262 26880 8558 26908
rect 8552 26868 8558 26880
rect 8610 26868 8616 26920
rect 8828 26868 8834 26920
rect 8886 26908 8892 26920
rect 20696 26908 20702 26920
rect 8886 26880 20702 26908
rect 8886 26868 8892 26880
rect 20696 26868 20702 26880
rect 20754 26868 20760 26920
rect 25940 26868 25946 26920
rect 25998 26908 26004 26920
rect 26124 26908 26130 26920
rect 25998 26880 26130 26908
rect 25998 26868 26004 26880
rect 26124 26868 26130 26880
rect 26182 26868 26188 26920
rect 37995 26911 38053 26917
rect 37995 26908 38007 26911
rect 26234 26880 38007 26908
rect 16556 26800 16562 26852
rect 16614 26840 16620 26852
rect 22996 26840 23002 26852
rect 16614 26812 23002 26840
rect 16614 26800 16620 26812
rect 22996 26800 23002 26812
rect 23054 26800 23060 26852
rect 24652 26800 24658 26852
rect 24710 26840 24716 26852
rect 26234 26840 26262 26880
rect 37995 26877 38007 26880
rect 38041 26877 38053 26911
rect 37995 26871 38053 26877
rect 24710 26812 26262 26840
rect 24710 26800 24716 26812
rect 7816 26732 7822 26784
rect 7874 26772 7880 26784
rect 8184 26772 8190 26784
rect 7874 26744 8190 26772
rect 7874 26732 7880 26744
rect 8184 26732 8190 26744
rect 8242 26732 8248 26784
rect 8690 26732 8696 26784
rect 8748 26732 8754 26784
rect 21711 26775 21769 26781
rect 21711 26741 21723 26775
rect 21757 26772 21769 26775
rect 29620 26772 29626 26784
rect 21757 26744 29626 26772
rect 21757 26741 21769 26744
rect 21711 26735 21769 26741
rect 29620 26732 29626 26744
rect 29678 26732 29684 26784
rect 1086 26682 58862 26704
rect 1086 26630 19588 26682
rect 19640 26630 19652 26682
rect 19704 26630 19716 26682
rect 19768 26630 19780 26682
rect 19832 26630 50308 26682
rect 50360 26630 50372 26682
rect 50424 26630 50436 26682
rect 50488 26630 50500 26682
rect 50552 26630 58862 26682
rect 1086 26608 58862 26630
rect 8690 26528 8696 26580
rect 8748 26568 8754 26580
rect 22904 26568 22910 26580
rect 8748 26540 22910 26568
rect 8748 26528 8754 26540
rect 22904 26528 22910 26540
rect 22962 26528 22968 26580
rect 6804 26392 6810 26444
rect 6862 26432 6868 26444
rect 43515 26435 43573 26441
rect 43515 26432 43527 26435
rect 6862 26404 43527 26432
rect 6862 26392 6868 26404
rect 43515 26401 43527 26404
rect 43561 26401 43573 26435
rect 43515 26395 43573 26401
rect 12140 26324 12146 26376
rect 12198 26364 12204 26376
rect 29163 26367 29221 26373
rect 29163 26364 29175 26367
rect 12198 26336 29175 26364
rect 12198 26324 12204 26336
rect 29163 26333 29175 26336
rect 29209 26333 29221 26367
rect 29163 26327 29221 26333
rect 32932 26324 32938 26376
rect 32990 26364 32996 26376
rect 49127 26367 49185 26373
rect 49127 26364 49139 26367
rect 32990 26336 49139 26364
rect 32990 26324 32996 26336
rect 49127 26333 49139 26336
rect 49173 26333 49185 26367
rect 49127 26327 49185 26333
rect 25020 26296 25026 26308
rect 24981 26268 25026 26296
rect 25020 26256 25026 26268
rect 25078 26256 25084 26308
rect 31644 26256 31650 26308
rect 31702 26296 31708 26308
rect 34131 26299 34189 26305
rect 34131 26296 34143 26299
rect 31702 26268 34143 26296
rect 31702 26256 31708 26268
rect 34131 26265 34143 26268
rect 34177 26265 34189 26299
rect 34131 26259 34189 26265
rect 38728 26188 38734 26240
rect 38786 26228 38792 26240
rect 39004 26228 39010 26240
rect 38786 26200 39010 26228
rect 38786 26188 38792 26200
rect 39004 26188 39010 26200
rect 39062 26188 39068 26240
rect 1086 26138 58862 26160
rect 1086 26086 4228 26138
rect 4280 26086 4292 26138
rect 4344 26086 4356 26138
rect 4408 26086 4420 26138
rect 4472 26086 34948 26138
rect 35000 26086 35012 26138
rect 35064 26086 35076 26138
rect 35128 26086 35140 26138
rect 35192 26086 58862 26138
rect 1086 26064 58862 26086
rect 13612 26024 13618 26036
rect 13573 25996 13618 26024
rect 13612 25984 13618 25996
rect 13670 25984 13676 26036
rect 10211 25891 10269 25897
rect 10211 25888 10223 25891
rect 10134 25860 10223 25888
rect 8552 25820 8558 25832
rect 8446 25792 8558 25820
rect 8552 25780 8558 25792
rect 8610 25780 8616 25832
rect 8248 25696 8276 25772
rect 10134 25752 10162 25860
rect 10211 25857 10223 25860
rect 10257 25857 10269 25891
rect 10211 25851 10269 25857
rect 20328 25848 20334 25900
rect 20386 25888 20392 25900
rect 20386 25860 27550 25888
rect 20386 25848 20392 25860
rect 27522 25820 27550 25860
rect 37624 25820 37630 25832
rect 27522 25792 37630 25820
rect 37624 25780 37630 25792
rect 37682 25780 37688 25832
rect 42227 25823 42285 25829
rect 42227 25789 42239 25823
rect 42273 25789 42285 25823
rect 42227 25783 42285 25789
rect 20328 25752 20334 25764
rect 10134 25724 20334 25752
rect 20328 25712 20334 25724
rect 20386 25712 20392 25764
rect 20420 25712 20426 25764
rect 20478 25752 20484 25764
rect 42242 25752 42270 25783
rect 20478 25724 42270 25752
rect 20478 25712 20484 25724
rect 8184 25644 8190 25696
rect 8242 25656 8276 25696
rect 8242 25644 8248 25656
rect 8690 25644 8696 25696
rect 8748 25644 8754 25696
rect 8828 25644 8834 25696
rect 8886 25684 8892 25696
rect 22444 25684 22450 25696
rect 8886 25656 22450 25684
rect 8886 25644 8892 25656
rect 22444 25644 22450 25656
rect 22502 25644 22508 25696
rect 1086 25594 58862 25616
rect 1086 25542 19588 25594
rect 19640 25542 19652 25594
rect 19704 25542 19716 25594
rect 19768 25542 19780 25594
rect 19832 25542 50308 25594
rect 50360 25542 50372 25594
rect 50424 25542 50436 25594
rect 50488 25542 50500 25594
rect 50552 25542 58862 25594
rect 1086 25520 58862 25542
rect 8184 25440 8190 25492
rect 8242 25480 8248 25492
rect 22628 25480 22634 25492
rect 8242 25452 22634 25480
rect 8242 25440 8248 25452
rect 22628 25440 22634 25452
rect 22686 25440 22692 25492
rect 8690 25372 8696 25424
rect 8748 25412 8754 25424
rect 21616 25412 21622 25424
rect 8748 25384 21622 25412
rect 8748 25372 8754 25384
rect 21616 25372 21622 25384
rect 21674 25372 21680 25424
rect 37624 25236 37630 25288
rect 37682 25276 37688 25288
rect 44800 25276 44806 25288
rect 37682 25248 44806 25276
rect 37682 25236 37688 25248
rect 44800 25236 44806 25248
rect 44858 25236 44864 25288
rect 31552 25100 31558 25152
rect 31610 25140 31616 25152
rect 51703 25143 51761 25149
rect 51703 25140 51715 25143
rect 31610 25112 51715 25140
rect 31610 25100 31616 25112
rect 51703 25109 51715 25112
rect 51749 25109 51761 25143
rect 51703 25103 51761 25109
rect 1086 25050 58862 25072
rect 1086 24998 4228 25050
rect 4280 24998 4292 25050
rect 4344 24998 4356 25050
rect 4408 24998 4420 25050
rect 4472 24998 34948 25050
rect 35000 24998 35012 25050
rect 35064 24998 35076 25050
rect 35128 24998 35140 25050
rect 35192 24998 58862 25050
rect 1086 24976 58862 24998
rect 2204 24896 2210 24948
rect 2262 24936 2268 24948
rect 2572 24936 2578 24948
rect 2262 24908 2578 24936
rect 2262 24896 2268 24908
rect 2572 24896 2578 24908
rect 2630 24896 2636 24948
rect 7632 24936 7638 24948
rect 7558 24908 7638 24936
rect 7558 24880 7586 24908
rect 7632 24896 7638 24908
rect 7690 24896 7696 24948
rect 7540 24828 7546 24880
rect 7598 24828 7604 24880
rect 8828 24862 8834 24914
rect 8886 24862 8892 24914
rect 9012 24896 9018 24948
rect 9070 24936 9076 24948
rect 21524 24936 21530 24948
rect 9070 24908 21530 24936
rect 9070 24896 9076 24908
rect 21524 24896 21530 24908
rect 21582 24896 21588 24948
rect 23272 24896 23278 24948
rect 23330 24936 23336 24948
rect 23456 24936 23462 24948
rect 23330 24908 23462 24936
rect 23330 24896 23336 24908
rect 23456 24896 23462 24908
rect 23514 24896 23520 24948
rect 45536 24828 45542 24880
rect 45594 24868 45600 24880
rect 45720 24868 45726 24880
rect 45594 24840 45726 24868
rect 45594 24828 45600 24840
rect 45720 24828 45726 24840
rect 45778 24828 45784 24880
rect 8923 24803 8981 24809
rect 2480 24732 2486 24744
rect 2441 24704 2486 24732
rect 2480 24692 2486 24704
rect 2538 24692 2544 24744
rect 8248 24596 8276 24786
rect 8923 24769 8935 24803
rect 8969 24800 8981 24803
rect 20880 24800 20886 24812
rect 8969 24772 20886 24800
rect 8969 24769 8981 24772
rect 8923 24763 8981 24769
rect 20880 24760 20886 24772
rect 20938 24760 20944 24812
rect 20972 24732 20978 24744
rect 8432 24676 8460 24718
rect 8432 24636 8466 24676
rect 8460 24624 8466 24636
rect 8518 24624 8524 24676
rect 8598 24658 8604 24710
rect 8656 24658 8662 24710
rect 8814 24704 20978 24732
rect 20972 24692 20978 24704
rect 21030 24692 21036 24744
rect 9012 24624 9018 24676
rect 9070 24664 9076 24676
rect 21708 24664 21714 24676
rect 9070 24636 21714 24664
rect 9070 24624 9076 24636
rect 21708 24624 21714 24636
rect 21766 24624 21772 24676
rect 8923 24599 8981 24605
rect 8923 24596 8935 24599
rect 8248 24568 8935 24596
rect 8923 24565 8935 24568
rect 8969 24565 8981 24599
rect 8923 24559 8981 24565
rect 1086 24506 58862 24528
rect 1086 24454 19588 24506
rect 19640 24454 19652 24506
rect 19704 24454 19716 24506
rect 19768 24454 19780 24506
rect 19832 24454 50308 24506
rect 50360 24454 50372 24506
rect 50424 24454 50436 24506
rect 50488 24454 50500 24506
rect 50552 24454 58862 24506
rect 1086 24432 58862 24454
rect 8460 24352 8466 24404
rect 8518 24392 8524 24404
rect 21800 24392 21806 24404
rect 8518 24364 21806 24392
rect 8518 24352 8524 24364
rect 21800 24352 21806 24364
rect 21858 24352 21864 24404
rect 2480 24284 2486 24336
rect 2538 24324 2544 24336
rect 28424 24324 28430 24336
rect 2538 24296 28430 24324
rect 2538 24284 2544 24296
rect 28424 24284 28430 24296
rect 28482 24284 28488 24336
rect 43604 24256 43610 24268
rect 43565 24228 43610 24256
rect 43604 24216 43610 24228
rect 43662 24216 43668 24268
rect 7632 24148 7638 24200
rect 7690 24188 7696 24200
rect 32104 24188 32110 24200
rect 7690 24160 32110 24188
rect 7690 24148 7696 24160
rect 32104 24148 32110 24160
rect 32162 24148 32168 24200
rect 56576 24148 56582 24200
rect 56634 24188 56640 24200
rect 56760 24188 56766 24200
rect 56634 24160 56766 24188
rect 56634 24148 56640 24160
rect 56760 24148 56766 24160
rect 56818 24148 56824 24200
rect 12784 24080 12790 24132
rect 12842 24120 12848 24132
rect 20328 24120 20334 24132
rect 12842 24092 20334 24120
rect 12842 24080 12848 24092
rect 20328 24080 20334 24092
rect 20386 24080 20392 24132
rect 6712 24012 6718 24064
rect 6770 24052 6776 24064
rect 28519 24055 28577 24061
rect 28519 24052 28531 24055
rect 6770 24024 28531 24052
rect 6770 24012 6776 24024
rect 28519 24021 28531 24024
rect 28565 24021 28577 24055
rect 28519 24015 28577 24021
rect 1086 23962 58862 23984
rect 1086 23910 4228 23962
rect 4280 23910 4292 23962
rect 4344 23910 4356 23962
rect 4408 23910 4420 23962
rect 4472 23910 34948 23962
rect 35000 23910 35012 23962
rect 35064 23910 35076 23962
rect 35128 23910 35140 23962
rect 35192 23910 58862 23962
rect 1086 23888 58862 23910
rect 7632 23848 7638 23860
rect 7593 23820 7638 23848
rect 7632 23808 7638 23820
rect 7690 23808 7696 23860
rect 8644 23808 8650 23860
rect 8702 23808 8708 23860
rect 8828 23808 8834 23860
rect 8886 23848 8892 23860
rect 18215 23851 18273 23857
rect 8886 23820 13014 23848
rect 8886 23808 8892 23820
rect 12876 23780 12882 23792
rect 12837 23752 12882 23780
rect 12876 23740 12882 23752
rect 12934 23740 12940 23792
rect 12986 23712 13014 23820
rect 18215 23817 18227 23851
rect 18261 23848 18273 23851
rect 27044 23848 27050 23860
rect 18261 23820 27050 23848
rect 18261 23817 18273 23820
rect 18215 23811 18273 23817
rect 27044 23808 27050 23820
rect 27102 23808 27108 23860
rect 13060 23740 13066 23792
rect 13118 23780 13124 23792
rect 19963 23783 20021 23789
rect 19963 23780 19975 23783
rect 13118 23752 19975 23780
rect 13118 23740 13124 23752
rect 19963 23749 19975 23752
rect 20009 23749 20021 23783
rect 19963 23743 20021 23749
rect 18764 23712 18770 23724
rect 8630 23684 12922 23712
rect 12986 23684 18770 23712
rect 12143 23647 12201 23653
rect 8248 23508 8276 23596
rect 8414 23570 8420 23622
rect 8472 23570 8478 23622
rect 12143 23613 12155 23647
rect 12189 23644 12201 23647
rect 12784 23644 12790 23656
rect 12189 23616 12790 23644
rect 12189 23613 12201 23616
rect 12143 23607 12201 23613
rect 12784 23604 12790 23616
rect 12842 23604 12848 23656
rect 12894 23644 12922 23684
rect 18764 23672 18770 23684
rect 18822 23672 18828 23724
rect 20144 23644 20150 23656
rect 12894 23616 20150 23644
rect 20144 23604 20150 23616
rect 20202 23604 20208 23656
rect 8736 23536 8742 23588
rect 8794 23576 8800 23588
rect 8794 23548 12830 23576
rect 8794 23536 8800 23548
rect 12143 23511 12201 23517
rect 12143 23508 12155 23511
rect 8248 23480 12155 23508
rect 12143 23477 12155 23480
rect 12189 23477 12201 23511
rect 12802 23508 12830 23548
rect 12876 23536 12882 23588
rect 12934 23576 12940 23588
rect 32472 23576 32478 23588
rect 12934 23548 32478 23576
rect 12934 23536 12940 23548
rect 32472 23536 32478 23548
rect 32530 23536 32536 23588
rect 20236 23508 20242 23520
rect 12802 23480 20242 23508
rect 12143 23471 12201 23477
rect 20236 23468 20242 23480
rect 20294 23468 20300 23520
rect 1086 23418 58862 23440
rect 1086 23366 19588 23418
rect 19640 23366 19652 23418
rect 19704 23366 19716 23418
rect 19768 23366 19780 23418
rect 19832 23366 50308 23418
rect 50360 23366 50372 23418
rect 50424 23366 50436 23418
rect 50488 23366 50500 23418
rect 50552 23366 58862 23418
rect 1086 23344 58862 23366
rect 26492 22924 26498 22976
rect 26550 22964 26556 22976
rect 26676 22964 26682 22976
rect 26550 22936 26682 22964
rect 26550 22924 26556 22936
rect 26676 22924 26682 22936
rect 26734 22924 26740 22976
rect 1086 22874 58862 22896
rect 1086 22822 4228 22874
rect 4280 22822 4292 22874
rect 4344 22822 4356 22874
rect 4408 22822 4420 22874
rect 4472 22822 34948 22874
rect 35000 22822 35012 22874
rect 35064 22822 35076 22874
rect 35128 22822 35140 22874
rect 35192 22822 58862 22874
rect 1086 22800 58862 22822
rect 9107 22763 9165 22769
rect 9107 22760 9119 22763
rect 8800 22732 9119 22760
rect 8800 22610 8828 22732
rect 9107 22729 9119 22732
rect 9153 22729 9165 22763
rect 18396 22760 18402 22772
rect 9274 22732 18402 22760
rect 9107 22723 9165 22729
rect 18396 22720 18402 22732
rect 18454 22720 18460 22772
rect 9291 22627 9349 22633
rect 9291 22624 9303 22627
rect 8998 22596 9058 22624
rect 9182 22596 9303 22624
rect 9030 22420 9058 22596
rect 9291 22593 9303 22596
rect 9337 22593 9349 22627
rect 9291 22587 9349 22593
rect 33024 22584 33030 22636
rect 33082 22624 33088 22636
rect 55935 22627 55993 22633
rect 55935 22624 55947 22627
rect 33082 22596 55947 22624
rect 33082 22584 33088 22596
rect 55935 22593 55947 22596
rect 55981 22593 55993 22627
rect 55935 22587 55993 22593
rect 9107 22559 9165 22565
rect 9107 22525 9119 22559
rect 9153 22556 9165 22559
rect 18304 22556 18310 22568
rect 9153 22528 18310 22556
rect 9153 22525 9165 22528
rect 9107 22519 9165 22525
rect 18304 22516 18310 22528
rect 18362 22516 18368 22568
rect 25940 22516 25946 22568
rect 25998 22556 26004 22568
rect 36155 22559 36213 22565
rect 36155 22556 36167 22559
rect 25998 22528 36167 22556
rect 25998 22516 26004 22528
rect 36155 22525 36167 22528
rect 36201 22525 36213 22559
rect 36155 22519 36213 22525
rect 9291 22491 9349 22497
rect 9291 22457 9303 22491
rect 9337 22488 9349 22491
rect 18028 22488 18034 22500
rect 9337 22460 18034 22488
rect 9337 22457 9349 22460
rect 9291 22451 9349 22457
rect 18028 22448 18034 22460
rect 18086 22448 18092 22500
rect 18488 22420 18494 22432
rect 9030 22392 18494 22420
rect 18488 22380 18494 22392
rect 18546 22380 18552 22432
rect 1086 22330 58862 22352
rect 1086 22278 19588 22330
rect 19640 22278 19652 22330
rect 19704 22278 19716 22330
rect 19768 22278 19780 22330
rect 19832 22278 50308 22330
rect 50360 22278 50372 22330
rect 50424 22278 50436 22330
rect 50488 22278 50500 22330
rect 50552 22278 58862 22330
rect 1086 22256 58862 22278
rect 2851 22151 2909 22157
rect 2851 22117 2863 22151
rect 2897 22148 2909 22151
rect 33760 22148 33766 22160
rect 2897 22120 33766 22148
rect 2897 22117 2909 22120
rect 2851 22111 2909 22117
rect 33760 22108 33766 22120
rect 33818 22108 33824 22160
rect 22002 21984 22122 22012
rect 17663 21947 17721 21953
rect 17663 21913 17675 21947
rect 17709 21944 17721 21947
rect 22002 21944 22030 21984
rect 17709 21916 22030 21944
rect 17709 21913 17721 21916
rect 17663 21907 17721 21913
rect 13428 21836 13434 21888
rect 13486 21876 13492 21888
rect 21067 21879 21125 21885
rect 21067 21876 21079 21879
rect 13486 21848 21079 21876
rect 13486 21836 13492 21848
rect 21067 21845 21079 21848
rect 21113 21845 21125 21879
rect 22094 21876 22122 21984
rect 46827 21947 46885 21953
rect 46827 21913 46839 21947
rect 46873 21944 46885 21947
rect 50596 21944 50602 21956
rect 46873 21916 50602 21944
rect 46873 21913 46885 21916
rect 46827 21907 46885 21913
rect 50596 21904 50602 21916
rect 50654 21904 50660 21956
rect 35508 21876 35514 21888
rect 22094 21848 35514 21876
rect 21067 21839 21125 21845
rect 35508 21836 35514 21848
rect 35566 21836 35572 21888
rect 47928 21876 47934 21888
rect 47889 21848 47934 21876
rect 47928 21836 47934 21848
rect 47986 21836 47992 21888
rect 1086 21786 58862 21808
rect 1086 21734 4228 21786
rect 4280 21734 4292 21786
rect 4344 21734 4356 21786
rect 4408 21734 4420 21786
rect 4472 21734 34948 21786
rect 35000 21734 35012 21786
rect 35064 21734 35076 21786
rect 35128 21734 35140 21786
rect 35192 21734 58862 21786
rect 1086 21712 58862 21734
rect 8555 21675 8613 21681
rect 8555 21672 8567 21675
rect 8248 21644 8567 21672
rect 8248 21556 8276 21644
rect 8555 21641 8567 21644
rect 8601 21641 8613 21675
rect 8555 21635 8613 21641
rect 17016 21536 17022 21548
rect 8446 21508 17022 21536
rect 17016 21496 17022 21508
rect 17074 21496 17080 21548
rect 8555 21471 8613 21477
rect 8555 21437 8567 21471
rect 8601 21468 8613 21471
rect 16924 21468 16930 21480
rect 8601 21440 16930 21468
rect 8601 21437 8613 21440
rect 8555 21431 8613 21437
rect 16924 21428 16930 21440
rect 16982 21428 16988 21480
rect 30359 21471 30417 21477
rect 30359 21437 30371 21471
rect 30405 21468 30417 21471
rect 42132 21468 42138 21480
rect 30405 21440 42138 21468
rect 30405 21437 30417 21440
rect 30359 21431 30417 21437
rect 42132 21428 42138 21440
rect 42190 21428 42196 21480
rect 8460 21292 8466 21344
rect 8518 21292 8524 21344
rect 8644 21292 8650 21344
rect 8702 21332 8708 21344
rect 16832 21332 16838 21344
rect 8702 21304 16838 21332
rect 8702 21292 8708 21304
rect 16832 21292 16838 21304
rect 16890 21292 16896 21344
rect 1086 21242 58862 21264
rect 1086 21190 19588 21242
rect 19640 21190 19652 21242
rect 19704 21190 19716 21242
rect 19768 21190 19780 21242
rect 19832 21190 50308 21242
rect 50360 21190 50372 21242
rect 50424 21190 50436 21242
rect 50488 21190 50500 21242
rect 50552 21190 58862 21242
rect 1086 21168 58862 21190
rect 18764 20816 18770 20868
rect 18822 20856 18828 20868
rect 19960 20856 19966 20868
rect 18822 20828 19966 20856
rect 18822 20816 18828 20828
rect 19960 20816 19966 20828
rect 20018 20816 20024 20868
rect 1086 20698 58862 20720
rect 1086 20646 4228 20698
rect 4280 20646 4292 20698
rect 4344 20646 4356 20698
rect 4408 20646 4420 20698
rect 4472 20646 34948 20698
rect 35000 20646 35012 20698
rect 35064 20646 35076 20698
rect 35128 20646 35140 20698
rect 35192 20646 58862 20698
rect 1086 20624 58862 20646
rect 8460 20544 8466 20596
rect 8518 20544 8524 20596
rect 48112 20544 48118 20596
rect 48170 20584 48176 20596
rect 56487 20587 56545 20593
rect 56487 20584 56499 20587
rect 48170 20556 56499 20584
rect 48170 20544 48176 20556
rect 56487 20553 56499 20556
rect 56533 20553 56545 20587
rect 56487 20547 56545 20553
rect 17770 20488 20006 20516
rect 9472 20408 9478 20460
rect 9530 20448 9536 20460
rect 17770 20448 17798 20488
rect 9530 20420 17798 20448
rect 9530 20408 9536 20420
rect 10852 20380 10858 20392
rect 8248 20244 8276 20332
rect 8414 20306 8420 20358
rect 8472 20306 8478 20358
rect 8630 20352 10714 20380
rect 10813 20352 10858 20380
rect 10686 20312 10714 20352
rect 10852 20340 10858 20352
rect 10910 20340 10916 20392
rect 19978 20380 20006 20488
rect 48112 20380 48118 20392
rect 19978 20352 48118 20380
rect 48112 20340 48118 20352
rect 48170 20340 48176 20392
rect 16188 20312 16194 20324
rect 10686 20284 16194 20312
rect 16188 20272 16194 20284
rect 16246 20272 16252 20324
rect 14532 20244 14538 20256
rect 8248 20216 14538 20244
rect 14532 20204 14538 20216
rect 14590 20204 14596 20256
rect 1086 20154 58862 20176
rect 1086 20102 19588 20154
rect 19640 20102 19652 20154
rect 19704 20102 19716 20154
rect 19768 20102 19780 20154
rect 19832 20102 50308 20154
rect 50360 20102 50372 20154
rect 50424 20102 50436 20154
rect 50488 20102 50500 20154
rect 50552 20102 58862 20154
rect 1086 20080 58862 20102
rect 8460 20000 8466 20052
rect 8518 20040 8524 20052
rect 16280 20040 16286 20052
rect 8518 20012 16286 20040
rect 8518 20000 8524 20012
rect 16280 20000 16286 20012
rect 16338 20000 16344 20052
rect 19150 19876 27458 19904
rect 5608 19796 5614 19848
rect 5666 19836 5672 19848
rect 19150 19836 19178 19876
rect 27320 19836 27326 19848
rect 5666 19808 19178 19836
rect 20438 19808 27326 19836
rect 5666 19796 5672 19808
rect 10944 19728 10950 19780
rect 11002 19768 11008 19780
rect 20438 19768 20466 19808
rect 27320 19796 27326 19808
rect 27378 19796 27384 19848
rect 27430 19836 27458 19876
rect 49032 19836 49038 19848
rect 27430 19808 49038 19836
rect 49032 19796 49038 19808
rect 49090 19796 49096 19848
rect 42227 19771 42285 19777
rect 42227 19768 42239 19771
rect 11002 19740 20466 19768
rect 27338 19740 42239 19768
rect 11002 19728 11008 19740
rect 26032 19660 26038 19712
rect 26090 19700 26096 19712
rect 27338 19700 27366 19740
rect 42227 19737 42239 19740
rect 42273 19737 42285 19771
rect 42227 19731 42285 19737
rect 26090 19672 27366 19700
rect 26090 19660 26096 19672
rect 27412 19660 27418 19712
rect 27470 19700 27476 19712
rect 40295 19703 40353 19709
rect 40295 19700 40307 19703
rect 27470 19672 40307 19700
rect 27470 19660 27476 19672
rect 40295 19669 40307 19672
rect 40341 19669 40353 19703
rect 40295 19663 40353 19669
rect 1086 19610 58862 19632
rect 1086 19558 4228 19610
rect 4280 19558 4292 19610
rect 4344 19558 4356 19610
rect 4408 19558 4420 19610
rect 4472 19558 34948 19610
rect 35000 19558 35012 19610
rect 35064 19558 35076 19610
rect 35128 19558 35140 19610
rect 35192 19558 58862 19610
rect 1086 19536 58862 19558
rect 5608 19496 5614 19508
rect 5569 19468 5614 19496
rect 5608 19456 5614 19468
rect 5666 19456 5672 19508
rect 8460 19456 8466 19508
rect 8518 19456 8524 19508
rect 21340 19428 21346 19440
rect 21174 19400 21346 19428
rect 21174 19304 21202 19400
rect 21340 19388 21346 19400
rect 21398 19388 21404 19440
rect 26952 19320 26958 19372
rect 27010 19320 27016 19372
rect 37900 19320 37906 19372
rect 37958 19360 37964 19372
rect 37992 19360 37998 19372
rect 37958 19332 37998 19360
rect 37958 19320 37964 19332
rect 37992 19320 37998 19332
rect 38050 19320 38056 19372
rect 51056 19320 51062 19372
rect 51114 19360 51120 19372
rect 51240 19360 51246 19372
rect 51114 19332 51246 19360
rect 51114 19320 51120 19332
rect 51240 19320 51246 19332
rect 51298 19320 51304 19372
rect 7264 19292 7270 19304
rect 7225 19264 7270 19292
rect 7264 19252 7270 19264
rect 7322 19252 7328 19304
rect 8248 19168 8276 19244
rect 8414 19218 8420 19270
rect 8472 19218 8478 19270
rect 21156 19252 21162 19304
rect 21214 19252 21220 19304
rect 26970 19292 26998 19320
rect 27044 19292 27050 19304
rect 26970 19264 27050 19292
rect 27044 19252 27050 19264
rect 27102 19252 27108 19304
rect 20696 19184 20702 19236
rect 20754 19224 20760 19236
rect 23180 19224 23186 19236
rect 20754 19196 23186 19224
rect 20754 19184 20760 19196
rect 23180 19184 23186 19196
rect 23238 19184 23244 19236
rect 8184 19116 8190 19168
rect 8242 19128 8276 19168
rect 8242 19116 8248 19128
rect 8920 19116 8926 19168
rect 8978 19156 8984 19168
rect 13060 19156 13066 19168
rect 8978 19128 13066 19156
rect 8978 19116 8984 19128
rect 13060 19116 13066 19128
rect 13118 19116 13124 19168
rect 1086 19066 58862 19088
rect 1086 19014 19588 19066
rect 19640 19014 19652 19066
rect 19704 19014 19716 19066
rect 19768 19014 19780 19066
rect 19832 19014 50308 19066
rect 50360 19014 50372 19066
rect 50424 19014 50436 19066
rect 50488 19014 50500 19066
rect 50552 19014 58862 19066
rect 1086 18992 58862 19014
rect 8460 18912 8466 18964
rect 8518 18952 8524 18964
rect 10392 18952 10398 18964
rect 8518 18924 10398 18952
rect 8518 18912 8524 18924
rect 10392 18912 10398 18924
rect 10450 18912 10456 18964
rect 8552 18844 8558 18896
rect 8610 18884 8616 18896
rect 16740 18884 16746 18896
rect 8610 18856 16746 18884
rect 8610 18844 8616 18856
rect 16740 18844 16746 18856
rect 16798 18844 16804 18896
rect 27596 18708 27602 18760
rect 27654 18748 27660 18760
rect 27780 18748 27786 18760
rect 27654 18720 27786 18748
rect 27654 18708 27660 18720
rect 27780 18708 27786 18720
rect 27838 18708 27844 18760
rect 7264 18640 7270 18692
rect 7322 18680 7328 18692
rect 17936 18680 17942 18692
rect 7322 18652 17942 18680
rect 7322 18640 7328 18652
rect 17936 18640 17942 18652
rect 17994 18640 18000 18692
rect 2388 18572 2394 18624
rect 2446 18612 2452 18624
rect 35143 18615 35201 18621
rect 35143 18612 35155 18615
rect 2446 18584 35155 18612
rect 2446 18572 2452 18584
rect 35143 18581 35155 18584
rect 35189 18581 35201 18615
rect 35143 18575 35201 18581
rect 44987 18615 45045 18621
rect 44987 18581 44999 18615
rect 45033 18612 45045 18615
rect 47468 18612 47474 18624
rect 45033 18584 47474 18612
rect 45033 18581 45045 18584
rect 44987 18575 45045 18581
rect 47468 18572 47474 18584
rect 47526 18572 47532 18624
rect 1086 18522 58862 18544
rect 1086 18470 4228 18522
rect 4280 18470 4292 18522
rect 4344 18470 4356 18522
rect 4408 18470 4420 18522
rect 4472 18470 34948 18522
rect 35000 18470 35012 18522
rect 35064 18470 35076 18522
rect 35128 18470 35140 18522
rect 35192 18470 58862 18522
rect 1086 18448 58862 18470
rect 2575 18411 2633 18417
rect 2575 18377 2587 18411
rect 2621 18408 2633 18411
rect 7264 18408 7270 18420
rect 2621 18380 7270 18408
rect 2621 18377 2633 18380
rect 2575 18371 2633 18377
rect 7264 18368 7270 18380
rect 7322 18368 7328 18420
rect 8828 18368 8834 18420
rect 8886 18368 8892 18420
rect 9012 18368 9018 18420
rect 9070 18408 9076 18420
rect 14164 18408 14170 18420
rect 9070 18380 14170 18408
rect 9070 18368 9076 18380
rect 14164 18368 14170 18380
rect 14222 18368 14228 18420
rect 8647 18275 8705 18281
rect 8647 18272 8659 18275
rect 8446 18244 8659 18272
rect 8647 18241 8659 18244
rect 8693 18241 8705 18275
rect 9107 18275 9165 18281
rect 8647 18235 8705 18241
rect 8754 18244 8814 18272
rect 8754 18213 8782 18244
rect 9107 18241 9119 18275
rect 9153 18272 9165 18275
rect 13612 18272 13618 18284
rect 9153 18244 13618 18272
rect 9153 18241 9165 18244
rect 9107 18235 9165 18241
rect 13612 18232 13618 18244
rect 13670 18232 13676 18284
rect 8739 18207 8797 18213
rect 8739 18173 8751 18207
rect 8785 18173 8797 18207
rect 11496 18204 11502 18216
rect 8998 18176 11502 18204
rect 8739 18167 8797 18173
rect 11496 18164 11502 18176
rect 11554 18164 11560 18216
rect 47103 18207 47161 18213
rect 47103 18173 47115 18207
rect 47149 18204 47161 18207
rect 51700 18204 51706 18216
rect 47149 18176 51706 18204
rect 47149 18173 47161 18176
rect 47103 18167 47161 18173
rect 51700 18164 51706 18176
rect 51758 18164 51764 18216
rect 54003 18207 54061 18213
rect 54003 18173 54015 18207
rect 54049 18173 54061 18207
rect 54003 18167 54061 18173
rect 33208 18096 33214 18148
rect 33266 18136 33272 18148
rect 40660 18136 40666 18148
rect 33266 18108 40666 18136
rect 33266 18096 33272 18108
rect 40660 18096 40666 18108
rect 40718 18096 40724 18148
rect 44156 18096 44162 18148
rect 44214 18136 44220 18148
rect 54018 18136 54046 18167
rect 44214 18108 54046 18136
rect 44214 18096 44220 18108
rect 9015 18071 9073 18077
rect 9015 18037 9027 18071
rect 9061 18068 9073 18071
rect 12784 18068 12790 18080
rect 9061 18040 12790 18068
rect 9061 18037 9073 18040
rect 9015 18031 9073 18037
rect 12784 18028 12790 18040
rect 12842 18028 12848 18080
rect 1086 17978 58862 18000
rect 1086 17926 19588 17978
rect 19640 17926 19652 17978
rect 19704 17926 19716 17978
rect 19768 17926 19780 17978
rect 19832 17926 50308 17978
rect 50360 17926 50372 17978
rect 50424 17926 50436 17978
rect 50488 17926 50500 17978
rect 50552 17926 58862 17978
rect 1086 17904 58862 17926
rect 23919 17867 23977 17873
rect 23919 17833 23931 17867
rect 23965 17864 23977 17867
rect 27964 17864 27970 17876
rect 23965 17836 27970 17864
rect 23965 17833 23977 17836
rect 23919 17827 23977 17833
rect 27964 17824 27970 17836
rect 28022 17824 28028 17876
rect 8828 17756 8834 17808
rect 8886 17796 8892 17808
rect 56760 17796 56766 17808
rect 8886 17768 56766 17796
rect 8886 17756 8892 17768
rect 56760 17756 56766 17768
rect 56818 17756 56824 17808
rect 8736 17688 8742 17740
rect 8794 17728 8800 17740
rect 55196 17728 55202 17740
rect 8794 17700 55202 17728
rect 8794 17688 8800 17700
rect 55196 17688 55202 17700
rect 55254 17688 55260 17740
rect 1192 17620 1198 17672
rect 1250 17660 1256 17672
rect 35419 17663 35477 17669
rect 35419 17660 35431 17663
rect 1250 17632 35431 17660
rect 1250 17620 1256 17632
rect 35419 17629 35431 17632
rect 35465 17629 35477 17663
rect 39280 17660 39286 17672
rect 35419 17623 35477 17629
rect 35526 17632 39286 17660
rect 27964 17552 27970 17604
rect 28022 17592 28028 17604
rect 35526 17592 35554 17632
rect 39280 17620 39286 17632
rect 39338 17620 39344 17672
rect 28022 17564 35554 17592
rect 36538 17564 38406 17592
rect 28022 17552 28028 17564
rect 9383 17527 9441 17533
rect 9383 17493 9395 17527
rect 9429 17524 9441 17527
rect 19316 17524 19322 17536
rect 9429 17496 19322 17524
rect 9429 17493 9441 17496
rect 9383 17487 9441 17493
rect 19316 17484 19322 17496
rect 19374 17484 19380 17536
rect 23919 17527 23977 17533
rect 23919 17493 23931 17527
rect 23965 17524 23977 17527
rect 24195 17527 24253 17533
rect 24195 17524 24207 17527
rect 23965 17496 24207 17524
rect 23965 17493 23977 17496
rect 23919 17487 23977 17493
rect 24195 17493 24207 17496
rect 24241 17493 24253 17527
rect 24195 17487 24253 17493
rect 24560 17484 24566 17536
rect 24618 17524 24624 17536
rect 36538 17524 36566 17564
rect 24618 17496 36566 17524
rect 38179 17527 38237 17533
rect 24618 17484 24624 17496
rect 38179 17493 38191 17527
rect 38225 17524 38237 17527
rect 38268 17524 38274 17536
rect 38225 17496 38274 17524
rect 38225 17493 38237 17496
rect 38179 17487 38237 17493
rect 38268 17484 38274 17496
rect 38326 17484 38332 17536
rect 38378 17524 38406 17564
rect 48756 17524 48762 17536
rect 38378 17496 48762 17524
rect 48756 17484 48762 17496
rect 48814 17484 48820 17536
rect 1086 17434 58862 17456
rect 1086 17382 4228 17434
rect 4280 17382 4292 17434
rect 4344 17382 4356 17434
rect 4408 17382 4420 17434
rect 4472 17382 34948 17434
rect 35000 17382 35012 17434
rect 35064 17382 35076 17434
rect 35128 17382 35140 17434
rect 35192 17382 58862 17434
rect 1086 17360 58862 17382
rect 8000 17280 8006 17332
rect 8058 17280 8064 17332
rect 8828 17320 8834 17332
rect 8800 17280 8834 17320
rect 8886 17280 8892 17332
rect 7816 17076 7822 17128
rect 7874 17116 7880 17128
rect 8018 17116 8046 17280
rect 8800 17204 8828 17280
rect 9196 17246 9202 17298
rect 9254 17246 9260 17298
rect 23364 17280 23370 17332
rect 23422 17320 23428 17332
rect 33116 17320 33122 17332
rect 23422 17292 33122 17320
rect 23422 17280 23428 17292
rect 33116 17280 33122 17292
rect 33174 17280 33180 17332
rect 8736 17116 8742 17128
rect 7874 17088 8046 17116
rect 8446 17088 8742 17116
rect 7874 17076 7880 17088
rect 8736 17076 8742 17088
rect 8794 17076 8800 17128
rect 24560 17076 24566 17128
rect 24618 17116 24624 17128
rect 24744 17116 24750 17128
rect 24618 17088 24750 17116
rect 24618 17076 24624 17088
rect 24744 17076 24750 17088
rect 24802 17076 24808 17128
rect 1086 16890 58862 16912
rect 1086 16838 19588 16890
rect 19640 16838 19652 16890
rect 19704 16838 19716 16890
rect 19768 16838 19780 16890
rect 19832 16838 50308 16890
rect 50360 16838 50372 16890
rect 50424 16838 50436 16890
rect 50488 16838 50500 16890
rect 50552 16838 58862 16890
rect 1086 16816 58862 16838
rect 8644 16396 8650 16448
rect 8702 16436 8708 16448
rect 51056 16436 51062 16448
rect 8702 16408 51062 16436
rect 8702 16396 8708 16408
rect 51056 16396 51062 16408
rect 51114 16396 51120 16448
rect 1086 16346 58862 16368
rect 1086 16294 4228 16346
rect 4280 16294 4292 16346
rect 4344 16294 4356 16346
rect 4408 16294 4420 16346
rect 4472 16294 34948 16346
rect 35000 16294 35012 16346
rect 35064 16294 35076 16346
rect 35128 16294 35140 16346
rect 35192 16294 58862 16346
rect 1086 16272 58862 16294
rect 8736 16192 8742 16244
rect 8794 16192 8800 16244
rect 34683 16235 34741 16241
rect 34683 16201 34695 16235
rect 34729 16232 34741 16235
rect 36520 16232 36526 16244
rect 34729 16204 36526 16232
rect 34729 16201 34741 16204
rect 34683 16195 34741 16201
rect 36520 16192 36526 16204
rect 36578 16192 36584 16244
rect 8644 16074 8650 16126
rect 8702 16074 8708 16126
rect 24928 16124 24934 16176
rect 24986 16164 24992 16176
rect 27783 16167 27841 16173
rect 27783 16164 27795 16167
rect 24986 16136 27795 16164
rect 24986 16124 24992 16136
rect 27783 16133 27795 16136
rect 27829 16133 27841 16167
rect 27783 16127 27841 16133
rect 24560 16056 24566 16108
rect 24618 16096 24624 16108
rect 27875 16099 27933 16105
rect 27875 16096 27887 16099
rect 24618 16068 27887 16096
rect 24618 16056 24624 16068
rect 27875 16065 27887 16068
rect 27921 16065 27933 16099
rect 27875 16059 27933 16065
rect 2943 16031 3001 16037
rect 2943 15997 2955 16031
rect 2989 16028 3001 16031
rect 3032 16028 3038 16040
rect 2989 16000 3038 16028
rect 2989 15997 3001 16000
rect 2943 15991 3001 15997
rect 3032 15988 3038 16000
rect 3090 15988 3096 16040
rect 15084 15988 15090 16040
rect 15142 16028 15148 16040
rect 32659 16031 32717 16037
rect 32659 16028 32671 16031
rect 15142 16000 32671 16028
rect 15142 15988 15148 16000
rect 32659 15997 32671 16000
rect 32705 15997 32717 16031
rect 34588 16028 34594 16040
rect 34549 16000 34594 16028
rect 32659 15991 32717 15997
rect 34588 15988 34594 16000
rect 34646 15988 34652 16040
rect 34772 15988 34778 16040
rect 34830 16028 34836 16040
rect 35051 16031 35109 16037
rect 35051 16028 35063 16031
rect 34830 16000 35063 16028
rect 34830 15988 34836 16000
rect 35051 15997 35063 16000
rect 35097 15997 35109 16031
rect 35051 15991 35109 15997
rect 24744 15920 24750 15972
rect 24802 15960 24808 15972
rect 24928 15960 24934 15972
rect 24802 15932 24934 15960
rect 24802 15920 24808 15932
rect 24928 15920 24934 15932
rect 24986 15920 24992 15972
rect 27783 15963 27841 15969
rect 27783 15929 27795 15963
rect 27829 15960 27841 15963
rect 34683 15963 34741 15969
rect 34683 15960 34695 15963
rect 27829 15932 34695 15960
rect 27829 15929 27841 15932
rect 27783 15923 27841 15929
rect 34683 15929 34695 15932
rect 34729 15929 34741 15963
rect 34683 15923 34741 15929
rect 8736 15852 8742 15904
rect 8794 15892 8800 15904
rect 15176 15892 15182 15904
rect 8794 15864 15182 15892
rect 8794 15852 8800 15864
rect 15176 15852 15182 15864
rect 15234 15852 15240 15904
rect 1086 15802 58862 15824
rect 1086 15750 19588 15802
rect 19640 15750 19652 15802
rect 19704 15750 19716 15802
rect 19768 15750 19780 15802
rect 19832 15750 50308 15802
rect 50360 15750 50372 15802
rect 50424 15750 50436 15802
rect 50488 15750 50500 15802
rect 50552 15750 58862 15802
rect 1086 15728 58862 15750
rect 26679 15419 26737 15425
rect 26679 15385 26691 15419
rect 26725 15416 26737 15419
rect 50688 15416 50694 15428
rect 26725 15388 50694 15416
rect 26725 15385 26737 15388
rect 26679 15379 26737 15385
rect 50688 15376 50694 15388
rect 50746 15376 50752 15428
rect 45352 15308 45358 15360
rect 45410 15348 45416 15360
rect 45536 15348 45542 15360
rect 45410 15320 45542 15348
rect 45410 15308 45416 15320
rect 45536 15308 45542 15320
rect 45594 15308 45600 15360
rect 48204 15308 48210 15360
rect 48262 15348 48268 15360
rect 55935 15351 55993 15357
rect 55935 15348 55947 15351
rect 48262 15320 55947 15348
rect 48262 15308 48268 15320
rect 55935 15317 55947 15320
rect 55981 15317 55993 15351
rect 55935 15311 55993 15317
rect 1086 15258 58862 15280
rect 1086 15206 4228 15258
rect 4280 15206 4292 15258
rect 4344 15206 4356 15258
rect 4408 15206 4420 15258
rect 4472 15206 34948 15258
rect 35000 15206 35012 15258
rect 35064 15206 35076 15258
rect 35128 15206 35140 15258
rect 35192 15206 58862 15258
rect 1086 15184 58862 15206
rect 8460 15104 8466 15156
rect 8518 15104 8524 15156
rect 8644 15104 8650 15156
rect 8702 15144 8708 15156
rect 35324 15144 35330 15156
rect 8702 15116 35330 15144
rect 8702 15104 8708 15116
rect 35324 15104 35330 15116
rect 35382 15104 35388 15156
rect 13063 15079 13121 15085
rect 13063 15045 13075 15079
rect 13109 15076 13121 15079
rect 13796 15076 13802 15088
rect 13109 15048 13802 15076
rect 13109 15045 13121 15048
rect 13063 15039 13121 15045
rect 13796 15036 13802 15048
rect 13854 15036 13860 15088
rect 15179 15079 15237 15085
rect 15179 15045 15191 15079
rect 15225 15076 15237 15079
rect 18672 15076 18678 15088
rect 15225 15048 18678 15076
rect 15225 15045 15237 15048
rect 15179 15039 15237 15045
rect 18672 15036 18678 15048
rect 18730 15036 18736 15088
rect 8644 14968 8650 15020
rect 8702 15008 8708 15020
rect 48388 15008 48394 15020
rect 8702 14980 48394 15008
rect 8702 14968 8708 14980
rect 48388 14968 48394 14980
rect 48446 14968 48452 15020
rect 2296 14900 2302 14952
rect 2354 14940 2360 14952
rect 4047 14943 4105 14949
rect 4047 14940 4059 14943
rect 2354 14912 4059 14940
rect 2354 14900 2360 14912
rect 4047 14909 4059 14912
rect 4093 14909 4105 14943
rect 4047 14903 4105 14909
rect 8368 14866 8374 14918
rect 8426 14866 8432 14918
rect 29620 14900 29626 14952
rect 29678 14940 29684 14952
rect 31187 14943 31245 14949
rect 31187 14940 31199 14943
rect 29678 14912 31199 14940
rect 29678 14900 29684 14912
rect 31187 14909 31199 14912
rect 31233 14909 31245 14943
rect 31187 14903 31245 14909
rect 46824 14900 46830 14952
rect 46882 14940 46888 14952
rect 57683 14943 57741 14949
rect 57683 14940 57695 14943
rect 46882 14912 57695 14940
rect 46882 14900 46888 14912
rect 57683 14909 57695 14912
rect 57729 14909 57741 14943
rect 57683 14903 57741 14909
rect 1086 14714 58862 14736
rect 1086 14662 19588 14714
rect 19640 14662 19652 14714
rect 19704 14662 19716 14714
rect 19768 14662 19780 14714
rect 19832 14662 50308 14714
rect 50360 14662 50372 14714
rect 50424 14662 50436 14714
rect 50488 14662 50500 14714
rect 50552 14662 58862 14714
rect 1086 14640 58862 14662
rect 18396 14492 18402 14544
rect 18454 14532 18460 14544
rect 18856 14532 18862 14544
rect 18454 14504 18862 14532
rect 18454 14492 18460 14504
rect 18856 14492 18862 14504
rect 18914 14492 18920 14544
rect 44616 14464 44622 14476
rect 44577 14436 44622 14464
rect 44616 14424 44622 14436
rect 44674 14424 44680 14476
rect 6988 14356 6994 14408
rect 7046 14396 7052 14408
rect 25664 14396 25670 14408
rect 7046 14368 25670 14396
rect 7046 14356 7052 14368
rect 25664 14356 25670 14368
rect 25722 14356 25728 14408
rect 7632 14288 7638 14340
rect 7690 14328 7696 14340
rect 30819 14331 30877 14337
rect 30819 14328 30831 14331
rect 7690 14300 30831 14328
rect 7690 14288 7696 14300
rect 30819 14297 30831 14300
rect 30865 14297 30877 14331
rect 30819 14291 30877 14297
rect 25756 14260 25762 14272
rect 25717 14232 25762 14260
rect 25756 14220 25762 14232
rect 25814 14220 25820 14272
rect 36983 14263 37041 14269
rect 36983 14229 36995 14263
rect 37029 14260 37041 14263
rect 45168 14260 45174 14272
rect 37029 14232 45174 14260
rect 37029 14229 37041 14232
rect 36983 14223 37041 14229
rect 45168 14220 45174 14232
rect 45226 14220 45232 14272
rect 52344 14220 52350 14272
rect 52402 14260 52408 14272
rect 52991 14263 53049 14269
rect 52991 14260 53003 14263
rect 52402 14232 53003 14260
rect 52402 14220 52408 14232
rect 52991 14229 53003 14232
rect 53037 14229 53049 14263
rect 52991 14223 53049 14229
rect 1086 14170 58862 14192
rect 1086 14118 4228 14170
rect 4280 14118 4292 14170
rect 4344 14118 4356 14170
rect 4408 14118 4420 14170
rect 4472 14118 34948 14170
rect 35000 14118 35012 14170
rect 35064 14118 35076 14170
rect 35128 14118 35140 14170
rect 35192 14118 58862 14170
rect 1086 14096 58862 14118
rect 6988 14056 6994 14068
rect 6949 14028 6994 14056
rect 6988 14016 6994 14028
rect 7046 14016 7052 14068
rect 10576 14016 10582 14068
rect 10634 14056 10640 14068
rect 25756 14056 25762 14068
rect 10634 14028 25762 14056
rect 10634 14016 10640 14028
rect 25756 14016 25762 14028
rect 25814 14016 25820 14068
rect 26035 13991 26093 13997
rect 26035 13957 26047 13991
rect 26081 13988 26093 13991
rect 40660 13988 40666 14000
rect 26081 13960 40666 13988
rect 26081 13957 26093 13960
rect 26035 13951 26093 13957
rect 40660 13948 40666 13960
rect 40718 13948 40724 14000
rect 32380 13920 32386 13932
rect 8354 13892 32386 13920
rect 32380 13880 32386 13892
rect 32438 13880 32444 13932
rect 8000 13812 8006 13864
rect 8058 13852 8064 13864
rect 8058 13824 8262 13852
rect 8058 13812 8064 13824
rect 12508 13812 12514 13864
rect 12566 13852 12572 13864
rect 45536 13852 45542 13864
rect 12566 13824 45542 13852
rect 12566 13812 12572 13824
rect 45536 13812 45542 13824
rect 45594 13812 45600 13864
rect 49860 13784 49866 13796
rect 49821 13756 49866 13784
rect 49860 13744 49866 13756
rect 49918 13744 49924 13796
rect 1086 13626 58862 13648
rect 1086 13574 19588 13626
rect 19640 13574 19652 13626
rect 19704 13574 19716 13626
rect 19768 13574 19780 13626
rect 19832 13574 50308 13626
rect 50360 13574 50372 13626
rect 50424 13574 50436 13626
rect 50488 13574 50500 13626
rect 50552 13574 58862 13626
rect 1086 13552 58862 13574
rect 3676 13132 3682 13184
rect 3734 13172 3740 13184
rect 17108 13172 17114 13184
rect 3734 13144 17114 13172
rect 3734 13132 3740 13144
rect 17108 13132 17114 13144
rect 17166 13132 17172 13184
rect 1086 13082 58862 13104
rect 1086 13030 4228 13082
rect 4280 13030 4292 13082
rect 4344 13030 4356 13082
rect 4408 13030 4420 13082
rect 4472 13030 34948 13082
rect 35000 13030 35012 13082
rect 35064 13030 35076 13082
rect 35128 13030 35140 13082
rect 35192 13030 58862 13082
rect 1086 13008 58862 13030
rect 8138 12928 8144 12980
rect 8196 12928 8202 12980
rect 17108 12928 17114 12980
rect 17166 12968 17172 12980
rect 27783 12971 27841 12977
rect 27783 12968 27795 12971
rect 17166 12940 27795 12968
rect 17166 12928 17172 12940
rect 27783 12937 27795 12940
rect 27829 12937 27841 12971
rect 44708 12968 44714 12980
rect 44669 12940 44714 12968
rect 27783 12931 27841 12937
rect 44708 12928 44714 12940
rect 44766 12928 44772 12980
rect 52899 12903 52957 12909
rect 52899 12900 52911 12903
rect 22278 12872 52911 12900
rect 21340 12832 21346 12844
rect 8262 12804 21346 12832
rect 21340 12792 21346 12804
rect 21398 12792 21404 12844
rect 21892 12792 21898 12844
rect 21950 12832 21956 12844
rect 22278 12832 22306 12872
rect 52899 12869 52911 12872
rect 52945 12869 52957 12903
rect 52899 12863 52957 12869
rect 21950 12804 22306 12832
rect 21950 12792 21956 12804
rect 10760 12724 10766 12776
rect 10818 12764 10824 12776
rect 22171 12767 22229 12773
rect 22171 12764 22183 12767
rect 10818 12736 22183 12764
rect 10818 12724 10824 12736
rect 22171 12733 22183 12736
rect 22217 12733 22229 12767
rect 23824 12764 23830 12776
rect 23785 12736 23830 12764
rect 22171 12727 22229 12733
rect 23824 12724 23830 12736
rect 23882 12724 23888 12776
rect 42868 12764 42874 12776
rect 33042 12736 42874 12764
rect 21340 12656 21346 12708
rect 21398 12696 21404 12708
rect 33042 12696 33070 12736
rect 42868 12724 42874 12736
rect 42926 12724 42932 12776
rect 45815 12767 45873 12773
rect 45815 12733 45827 12767
rect 45861 12764 45873 12767
rect 51792 12764 51798 12776
rect 45861 12736 51798 12764
rect 45861 12733 45873 12736
rect 45815 12727 45873 12733
rect 51792 12724 51798 12736
rect 51850 12724 51856 12776
rect 21398 12668 33070 12696
rect 21398 12656 21404 12668
rect 1086 12538 58862 12560
rect 1086 12486 19588 12538
rect 19640 12486 19652 12538
rect 19704 12486 19716 12538
rect 19768 12486 19780 12538
rect 19832 12486 50308 12538
rect 50360 12486 50372 12538
rect 50424 12486 50436 12538
rect 50488 12486 50500 12538
rect 50552 12486 58862 12538
rect 1086 12464 58862 12486
rect 20331 12427 20389 12433
rect 20331 12393 20343 12427
rect 20377 12424 20389 12427
rect 21064 12424 21070 12436
rect 20377 12396 21070 12424
rect 20377 12393 20389 12396
rect 20331 12387 20389 12393
rect 21064 12384 21070 12396
rect 21122 12384 21128 12436
rect 11496 12316 11502 12368
rect 11554 12356 11560 12368
rect 13244 12356 13250 12368
rect 11554 12328 13250 12356
rect 11554 12316 11560 12328
rect 13244 12316 13250 12328
rect 13302 12316 13308 12368
rect 38470 12328 38682 12356
rect 7816 12248 7822 12300
rect 7874 12288 7880 12300
rect 24379 12291 24437 12297
rect 24379 12288 24391 12291
rect 7874 12260 24391 12288
rect 7874 12248 7880 12260
rect 24379 12257 24391 12260
rect 24425 12257 24437 12291
rect 24379 12251 24437 12257
rect 26216 12248 26222 12300
rect 26274 12288 26280 12300
rect 38470 12288 38498 12328
rect 26274 12260 38498 12288
rect 38654 12288 38682 12328
rect 48756 12316 48762 12368
rect 48814 12356 48820 12368
rect 49216 12356 49222 12368
rect 48814 12328 49222 12356
rect 48814 12316 48820 12328
rect 49216 12316 49222 12328
rect 49274 12316 49280 12368
rect 42227 12291 42285 12297
rect 42227 12288 42239 12291
rect 38654 12260 42239 12288
rect 26274 12248 26280 12260
rect 42227 12257 42239 12260
rect 42273 12257 42285 12291
rect 42227 12251 42285 12257
rect 6436 12180 6442 12232
rect 6494 12220 6500 12232
rect 6804 12220 6810 12232
rect 6494 12192 6810 12220
rect 6494 12180 6500 12192
rect 6804 12180 6810 12192
rect 6862 12180 6868 12232
rect 26216 12152 26222 12164
rect 11330 12124 26222 12152
rect 6804 12044 6810 12096
rect 6862 12084 6868 12096
rect 11330 12084 11358 12124
rect 26216 12112 26222 12124
rect 26274 12112 26280 12164
rect 6862 12056 11358 12084
rect 33303 12087 33361 12093
rect 6862 12044 6868 12056
rect 33303 12053 33315 12087
rect 33349 12084 33361 12087
rect 40292 12084 40298 12096
rect 33349 12056 40298 12084
rect 33349 12053 33361 12056
rect 33303 12047 33361 12053
rect 40292 12044 40298 12056
rect 40350 12044 40356 12096
rect 44064 12044 44070 12096
rect 44122 12084 44128 12096
rect 44435 12087 44493 12093
rect 44435 12084 44447 12087
rect 44122 12056 44447 12084
rect 44122 12044 44128 12056
rect 44435 12053 44447 12056
rect 44481 12053 44493 12087
rect 44435 12047 44493 12053
rect 1086 11994 58862 12016
rect 1086 11942 4228 11994
rect 4280 11942 4292 11994
rect 4344 11942 4356 11994
rect 4408 11942 4420 11994
rect 4472 11942 34948 11994
rect 35000 11942 35012 11994
rect 35064 11942 35076 11994
rect 35128 11942 35140 11994
rect 35192 11942 58862 11994
rect 1086 11920 58862 11942
rect 11680 11840 11686 11892
rect 11738 11880 11744 11892
rect 15176 11880 15182 11892
rect 11738 11852 15182 11880
rect 11738 11840 11744 11852
rect 15176 11840 15182 11852
rect 15234 11840 15240 11892
rect 6436 11704 6442 11756
rect 6494 11744 6500 11756
rect 6804 11744 6810 11756
rect 6494 11716 6810 11744
rect 6494 11704 6500 11716
rect 6804 11704 6810 11716
rect 6862 11704 6868 11756
rect 8092 11704 8098 11756
rect 8150 11744 8156 11756
rect 8150 11716 8262 11744
rect 8150 11704 8156 11716
rect 26216 11704 26222 11756
rect 26274 11744 26280 11756
rect 37348 11744 37354 11756
rect 26274 11716 37354 11744
rect 26274 11704 26280 11716
rect 37348 11704 37354 11716
rect 37406 11704 37412 11756
rect 19040 11676 19046 11688
rect 19001 11648 19046 11676
rect 19040 11636 19046 11648
rect 19098 11636 19104 11688
rect 49403 11679 49461 11685
rect 49403 11645 49415 11679
rect 49449 11645 49461 11679
rect 49403 11639 49461 11645
rect 55935 11679 55993 11685
rect 55935 11645 55947 11679
rect 55981 11676 55993 11679
rect 59704 11676 59710 11688
rect 55981 11648 59710 11676
rect 55981 11645 55993 11648
rect 55935 11639 55993 11645
rect 24836 11568 24842 11620
rect 24894 11608 24900 11620
rect 26216 11608 26222 11620
rect 24894 11580 26222 11608
rect 24894 11568 24900 11580
rect 26216 11568 26222 11580
rect 26274 11568 26280 11620
rect 37900 11540 37906 11552
rect 8354 11512 37906 11540
rect 37900 11500 37906 11512
rect 37958 11500 37964 11552
rect 49418 11540 49446 11639
rect 59704 11636 59710 11648
rect 59762 11636 59768 11688
rect 58600 11608 58606 11620
rect 53650 11580 58606 11608
rect 53650 11540 53678 11580
rect 58600 11568 58606 11580
rect 58658 11568 58664 11620
rect 49418 11512 53678 11540
rect 1086 11450 58862 11472
rect 1086 11398 19588 11450
rect 19640 11398 19652 11450
rect 19704 11398 19716 11450
rect 19768 11398 19780 11450
rect 19832 11398 50308 11450
rect 50360 11398 50372 11450
rect 50424 11398 50436 11450
rect 50488 11398 50500 11450
rect 50552 11398 58862 11450
rect 1086 11376 58862 11398
rect 9288 10956 9294 11008
rect 9346 10996 9352 11008
rect 33300 10996 33306 11008
rect 9346 10968 33306 10996
rect 9346 10956 9352 10968
rect 33300 10956 33306 10968
rect 33358 10956 33364 11008
rect 1086 10906 58862 10928
rect 1086 10854 4228 10906
rect 4280 10854 4292 10906
rect 4344 10854 4356 10906
rect 4408 10854 4420 10906
rect 4472 10854 34948 10906
rect 35000 10854 35012 10906
rect 35064 10854 35076 10906
rect 35128 10854 35140 10906
rect 35192 10854 58862 10906
rect 1086 10832 58862 10854
rect 8524 10764 19914 10792
rect 8524 10588 8552 10764
rect 19886 10656 19914 10764
rect 24836 10752 24842 10804
rect 24894 10792 24900 10804
rect 26216 10792 26222 10804
rect 24894 10764 26222 10792
rect 24894 10752 24900 10764
rect 26216 10752 26222 10764
rect 26274 10752 26280 10804
rect 29804 10792 29810 10804
rect 29765 10764 29810 10792
rect 29804 10752 29810 10764
rect 29862 10752 29868 10804
rect 19886 10628 20834 10656
rect 9656 10588 9662 10600
rect 8294 10560 8552 10588
rect 9550 10560 9662 10588
rect 8294 10472 8322 10560
rect 9656 10548 9662 10560
rect 9714 10548 9720 10600
rect 9840 10588 9846 10600
rect 9812 10548 9846 10588
rect 9898 10548 9904 10600
rect 20806 10588 20834 10628
rect 26216 10616 26222 10668
rect 26274 10656 26280 10668
rect 38636 10656 38642 10668
rect 26274 10628 38642 10656
rect 26274 10616 26280 10628
rect 38636 10616 38642 10628
rect 38694 10616 38700 10668
rect 24744 10588 24750 10600
rect 20806 10560 24750 10588
rect 24744 10548 24750 10560
rect 24802 10548 24808 10600
rect 9288 10480 9294 10532
rect 9346 10480 9352 10532
rect 9812 10472 9840 10548
rect 1086 10362 58862 10384
rect 1086 10310 19588 10362
rect 19640 10310 19652 10362
rect 19704 10310 19716 10362
rect 19768 10310 19780 10362
rect 19832 10310 50308 10362
rect 50360 10310 50372 10362
rect 50424 10310 50436 10362
rect 50488 10310 50500 10362
rect 50552 10310 58862 10362
rect 1086 10288 58862 10310
rect 9656 10208 9662 10260
rect 9714 10248 9720 10260
rect 34496 10248 34502 10260
rect 9714 10220 34502 10248
rect 9714 10208 9720 10220
rect 34496 10208 34502 10220
rect 34554 10208 34560 10260
rect 21340 10072 21346 10124
rect 21398 10112 21404 10124
rect 24008 10112 24014 10124
rect 21398 10084 24014 10112
rect 21398 10072 21404 10084
rect 24008 10072 24014 10084
rect 24066 10072 24072 10124
rect 2204 10004 2210 10056
rect 2262 10044 2268 10056
rect 32567 10047 32625 10053
rect 32567 10044 32579 10047
rect 2262 10016 32579 10044
rect 2262 10004 2268 10016
rect 32567 10013 32579 10016
rect 32613 10013 32625 10047
rect 32567 10007 32625 10013
rect 10392 9936 10398 9988
rect 10450 9976 10456 9988
rect 10668 9976 10674 9988
rect 10450 9948 10674 9976
rect 10450 9936 10456 9948
rect 10668 9936 10674 9948
rect 10726 9936 10732 9988
rect 24008 9936 24014 9988
rect 24066 9976 24072 9988
rect 33763 9979 33821 9985
rect 33763 9976 33775 9979
rect 24066 9948 33775 9976
rect 24066 9936 24072 9948
rect 33763 9945 33775 9948
rect 33809 9945 33821 9979
rect 33763 9939 33821 9945
rect 3860 9868 3866 9920
rect 3918 9908 3924 9920
rect 21340 9908 21346 9920
rect 3918 9880 21346 9908
rect 3918 9868 3924 9880
rect 21340 9868 21346 9880
rect 21398 9868 21404 9920
rect 32288 9908 32294 9920
rect 32249 9880 32294 9908
rect 32288 9868 32294 9880
rect 32346 9868 32352 9920
rect 49127 9911 49185 9917
rect 49127 9877 49139 9911
rect 49173 9908 49185 9911
rect 50136 9908 50142 9920
rect 49173 9880 50142 9908
rect 49173 9877 49185 9880
rect 49127 9871 49185 9877
rect 50136 9868 50142 9880
rect 50194 9868 50200 9920
rect 1086 9818 58862 9840
rect 1086 9766 4228 9818
rect 4280 9766 4292 9818
rect 4344 9766 4356 9818
rect 4408 9766 4420 9818
rect 4472 9766 34948 9818
rect 35000 9766 35012 9818
rect 35064 9766 35076 9818
rect 35128 9766 35140 9818
rect 35192 9766 58862 9818
rect 1086 9744 58862 9766
rect 6160 9704 6166 9716
rect 6086 9676 6166 9704
rect 6086 9648 6114 9676
rect 6160 9664 6166 9676
rect 6218 9664 6224 9716
rect 17476 9664 17482 9716
rect 17534 9704 17540 9716
rect 32288 9704 32294 9716
rect 17534 9676 32294 9704
rect 17534 9664 17540 9676
rect 32288 9664 32294 9676
rect 32346 9664 32352 9716
rect 41120 9664 41126 9716
rect 41178 9704 41184 9716
rect 44156 9704 44162 9716
rect 41178 9676 44162 9704
rect 41178 9664 41184 9676
rect 44156 9664 44162 9676
rect 44214 9664 44220 9716
rect 6068 9596 6074 9648
rect 6126 9596 6132 9648
rect 7724 9596 7730 9648
rect 7782 9636 7788 9648
rect 8092 9636 8098 9648
rect 7782 9608 8098 9636
rect 7782 9596 7788 9608
rect 8092 9596 8098 9608
rect 8150 9596 8156 9648
rect 10852 9596 10858 9648
rect 10910 9636 10916 9648
rect 11864 9636 11870 9648
rect 10910 9608 11870 9636
rect 10910 9596 10916 9608
rect 11864 9596 11870 9608
rect 11922 9596 11928 9648
rect 7540 9460 7546 9512
rect 7598 9500 7604 9512
rect 7724 9500 7730 9512
rect 7598 9472 7730 9500
rect 7598 9460 7604 9472
rect 7724 9460 7730 9472
rect 7782 9460 7788 9512
rect 10027 9503 10085 9509
rect 8368 9426 8374 9478
rect 8426 9426 8432 9478
rect 10027 9469 10039 9503
rect 10073 9500 10085 9503
rect 10852 9500 10858 9512
rect 10073 9472 10858 9500
rect 10073 9469 10085 9472
rect 10027 9463 10085 9469
rect 10852 9460 10858 9472
rect 10910 9460 10916 9512
rect 11036 9460 11042 9512
rect 11094 9500 11100 9512
rect 20791 9503 20849 9509
rect 20791 9500 20803 9503
rect 11094 9472 20803 9500
rect 11094 9460 11100 9472
rect 20791 9469 20803 9472
rect 20837 9469 20849 9503
rect 20791 9463 20849 9469
rect 31000 9432 31006 9444
rect 9490 9404 31006 9432
rect 9490 9384 9518 9404
rect 31000 9392 31006 9404
rect 31058 9392 31064 9444
rect 1086 9274 58862 9296
rect 1086 9222 19588 9274
rect 19640 9222 19652 9274
rect 19704 9222 19716 9274
rect 19768 9222 19780 9274
rect 19832 9222 50308 9274
rect 50360 9222 50372 9274
rect 50424 9222 50436 9274
rect 50488 9222 50500 9274
rect 50552 9222 58862 9274
rect 1086 9200 58862 9222
rect 8368 9120 8374 9172
rect 8426 9160 8432 9172
rect 29344 9160 29350 9172
rect 8426 9132 29350 9160
rect 8426 9120 8432 9132
rect 29344 9120 29350 9132
rect 29402 9120 29408 9172
rect 2848 8780 2854 8832
rect 2906 8820 2912 8832
rect 48388 8820 48394 8832
rect 2906 8792 48394 8820
rect 2906 8780 2912 8792
rect 48388 8780 48394 8792
rect 48446 8780 48452 8832
rect 1086 8730 58862 8752
rect 1086 8678 4228 8730
rect 4280 8678 4292 8730
rect 4344 8678 4356 8730
rect 4408 8678 4420 8730
rect 4472 8678 34948 8730
rect 35000 8678 35012 8730
rect 35064 8678 35076 8730
rect 35128 8678 35140 8730
rect 35192 8678 58862 8730
rect 1086 8656 58862 8678
rect 24008 8576 24014 8628
rect 24066 8616 24072 8628
rect 24066 8588 26814 8616
rect 24066 8576 24072 8588
rect 12235 8551 12293 8557
rect 12235 8517 12247 8551
rect 12281 8548 12293 8551
rect 26786 8548 26814 8588
rect 26952 8576 26958 8628
rect 27010 8616 27016 8628
rect 28240 8616 28246 8628
rect 27010 8588 28246 8616
rect 27010 8576 27016 8588
rect 28240 8576 28246 8588
rect 28298 8576 28304 8628
rect 48388 8616 48394 8628
rect 48349 8588 48394 8616
rect 48388 8576 48394 8588
rect 48446 8576 48452 8628
rect 39835 8551 39893 8557
rect 39835 8548 39847 8551
rect 12281 8520 26722 8548
rect 26786 8520 33070 8548
rect 12281 8517 12293 8520
rect 12235 8511 12293 8517
rect 3952 8480 3958 8492
rect 3913 8452 3958 8480
rect 3952 8440 3958 8452
rect 4010 8440 4016 8492
rect 8828 8440 8834 8492
rect 8886 8480 8892 8492
rect 26584 8480 26590 8492
rect 8886 8452 26590 8480
rect 8886 8440 8892 8452
rect 26584 8440 26590 8452
rect 26642 8440 26648 8492
rect 26694 8480 26722 8520
rect 26952 8480 26958 8492
rect 26694 8452 26958 8480
rect 26952 8440 26958 8452
rect 27010 8440 27016 8492
rect 33042 8480 33070 8520
rect 38654 8520 39847 8548
rect 38654 8480 38682 8520
rect 39835 8517 39847 8520
rect 39881 8517 39893 8551
rect 39835 8511 39893 8517
rect 40660 8508 40666 8560
rect 40718 8548 40724 8560
rect 41396 8548 41402 8560
rect 40718 8520 41402 8548
rect 40718 8508 40724 8520
rect 41396 8508 41402 8520
rect 41454 8508 41460 8560
rect 33042 8452 38682 8480
rect 8552 8412 8558 8424
rect 8262 8384 8558 8412
rect 8552 8372 8558 8384
rect 8610 8372 8616 8424
rect 12235 8415 12293 8421
rect 12235 8412 12247 8415
rect 10870 8384 12247 8412
rect 10870 8344 10898 8384
rect 12235 8381 12247 8384
rect 12281 8381 12293 8415
rect 12235 8375 12293 8381
rect 20696 8372 20702 8424
rect 20754 8412 20760 8424
rect 21432 8412 21438 8424
rect 20754 8384 21438 8412
rect 20754 8372 20760 8384
rect 21432 8372 21438 8384
rect 21490 8372 21496 8424
rect 47103 8415 47161 8421
rect 47103 8412 47115 8415
rect 22554 8384 47115 8412
rect 8570 8316 10898 8344
rect 8570 8296 8598 8316
rect 10944 8304 10950 8356
rect 11002 8344 11008 8356
rect 22554 8344 22582 8384
rect 47103 8381 47115 8384
rect 47149 8381 47161 8415
rect 47103 8375 47161 8381
rect 11002 8316 22582 8344
rect 11002 8304 11008 8316
rect 40292 8236 40298 8288
rect 40350 8276 40356 8288
rect 47284 8276 47290 8288
rect 40350 8248 47290 8276
rect 40350 8236 40356 8248
rect 47284 8236 47290 8248
rect 47342 8236 47348 8288
rect 1086 8186 58862 8208
rect 1086 8134 19588 8186
rect 19640 8134 19652 8186
rect 19704 8134 19716 8186
rect 19768 8134 19780 8186
rect 19832 8134 50308 8186
rect 50360 8134 50372 8186
rect 50424 8134 50436 8186
rect 50488 8134 50500 8186
rect 50552 8134 58862 8186
rect 1086 8112 58862 8134
rect 21064 8032 21070 8084
rect 21122 8072 21128 8084
rect 21616 8072 21622 8084
rect 21122 8044 21622 8072
rect 21122 8032 21128 8044
rect 21616 8032 21622 8044
rect 21674 8032 21680 8084
rect 22812 7896 22818 7948
rect 22870 7936 22876 7948
rect 23364 7936 23370 7948
rect 22870 7908 23370 7936
rect 22870 7896 22876 7908
rect 23364 7896 23370 7908
rect 23422 7896 23428 7948
rect 15636 7828 15642 7880
rect 15694 7868 15700 7880
rect 16372 7868 16378 7880
rect 15694 7840 16378 7868
rect 15694 7828 15700 7840
rect 16372 7828 16378 7840
rect 16430 7828 16436 7880
rect 22352 7828 22358 7880
rect 22410 7868 22416 7880
rect 22720 7868 22726 7880
rect 22410 7840 22726 7868
rect 22410 7828 22416 7840
rect 22720 7828 22726 7840
rect 22778 7828 22784 7880
rect 12232 7760 12238 7812
rect 12290 7800 12296 7812
rect 49311 7803 49369 7809
rect 49311 7800 49323 7803
rect 12290 7772 49323 7800
rect 12290 7760 12296 7772
rect 49311 7769 49323 7772
rect 49357 7769 49369 7803
rect 49311 7763 49369 7769
rect 15912 7692 15918 7744
rect 15970 7732 15976 7744
rect 16372 7732 16378 7744
rect 15970 7704 16378 7732
rect 15970 7692 15976 7704
rect 16372 7692 16378 7704
rect 16430 7692 16436 7744
rect 21340 7692 21346 7744
rect 21398 7732 21404 7744
rect 21800 7732 21806 7744
rect 21398 7704 21806 7732
rect 21398 7692 21404 7704
rect 21800 7692 21806 7704
rect 21858 7692 21864 7744
rect 22628 7692 22634 7744
rect 22686 7732 22692 7744
rect 22904 7732 22910 7744
rect 22686 7704 22910 7732
rect 22686 7692 22692 7704
rect 22904 7692 22910 7704
rect 22962 7692 22968 7744
rect 25112 7732 25118 7744
rect 25073 7704 25118 7732
rect 25112 7692 25118 7704
rect 25170 7692 25176 7744
rect 25572 7692 25578 7744
rect 25630 7732 25636 7744
rect 25940 7732 25946 7744
rect 25630 7704 25946 7732
rect 25630 7692 25636 7704
rect 25940 7692 25946 7704
rect 25998 7692 26004 7744
rect 46272 7732 46278 7744
rect 46233 7704 46278 7732
rect 46272 7692 46278 7704
rect 46330 7692 46336 7744
rect 1086 7642 58862 7664
rect 1086 7590 4228 7642
rect 4280 7590 4292 7642
rect 4344 7590 4356 7642
rect 4408 7590 4420 7642
rect 4472 7590 34948 7642
rect 35000 7590 35012 7642
rect 35064 7590 35076 7642
rect 35128 7590 35140 7642
rect 35192 7590 58862 7642
rect 1086 7568 58862 7590
rect 15820 7488 15826 7540
rect 15878 7528 15884 7540
rect 16280 7528 16286 7540
rect 15878 7500 16286 7528
rect 15878 7488 15884 7500
rect 16280 7488 16286 7500
rect 16338 7488 16344 7540
rect 18304 7488 18310 7540
rect 18362 7528 18368 7540
rect 18764 7528 18770 7540
rect 18362 7500 18770 7528
rect 18362 7488 18368 7500
rect 18764 7488 18770 7500
rect 18822 7488 18828 7540
rect 19408 7488 19414 7540
rect 19466 7528 19472 7540
rect 20328 7528 20334 7540
rect 19466 7500 20334 7528
rect 19466 7488 19472 7500
rect 20328 7488 20334 7500
rect 20386 7488 20392 7540
rect 22996 7488 23002 7540
rect 23054 7528 23060 7540
rect 23272 7528 23278 7540
rect 23054 7500 23278 7528
rect 23054 7488 23060 7500
rect 23272 7488 23278 7500
rect 23330 7488 23336 7540
rect 28976 7488 28982 7540
rect 29034 7528 29040 7540
rect 29988 7528 29994 7540
rect 29034 7500 29994 7528
rect 29034 7488 29040 7500
rect 29988 7488 29994 7500
rect 30046 7488 30052 7540
rect 31000 7488 31006 7540
rect 31058 7528 31064 7540
rect 46272 7528 46278 7540
rect 31058 7500 46278 7528
rect 31058 7488 31064 7500
rect 46272 7488 46278 7500
rect 46330 7488 46336 7540
rect 25112 7420 25118 7472
rect 25170 7460 25176 7472
rect 34680 7460 34686 7472
rect 25170 7432 34686 7460
rect 25170 7420 25176 7432
rect 34680 7420 34686 7432
rect 34738 7420 34744 7472
rect 8644 7352 8650 7404
rect 8702 7392 8708 7404
rect 23456 7392 23462 7404
rect 8702 7364 23462 7392
rect 8702 7352 8708 7364
rect 23456 7352 23462 7364
rect 23514 7352 23520 7404
rect 8368 7324 8374 7336
rect 8262 7296 8374 7324
rect 8368 7284 8374 7296
rect 8426 7284 8432 7336
rect 13983 7327 14041 7333
rect 13983 7293 13995 7327
rect 14029 7324 14041 7327
rect 16280 7324 16286 7336
rect 14029 7296 16286 7324
rect 14029 7293 14041 7296
rect 13983 7287 14041 7293
rect 16280 7284 16286 7296
rect 16338 7284 16344 7336
rect 24100 7188 24106 7200
rect 8538 7160 24106 7188
rect 24100 7148 24106 7160
rect 24158 7148 24164 7200
rect 1086 7098 58862 7120
rect 1086 7046 19588 7098
rect 19640 7046 19652 7098
rect 19704 7046 19716 7098
rect 19768 7046 19780 7098
rect 19832 7046 50308 7098
rect 50360 7046 50372 7098
rect 50424 7046 50436 7098
rect 50488 7046 50500 7098
rect 50552 7046 58862 7098
rect 1086 7024 58862 7046
rect 8184 6672 8190 6724
rect 8242 6712 8248 6724
rect 10024 6712 10030 6724
rect 8242 6684 10030 6712
rect 8242 6672 8248 6684
rect 10024 6672 10030 6684
rect 10082 6672 10088 6724
rect 5332 6604 5338 6656
rect 5390 6644 5396 6656
rect 5427 6647 5485 6653
rect 5427 6644 5439 6647
rect 5390 6616 5439 6644
rect 5390 6604 5396 6616
rect 5427 6613 5439 6616
rect 5473 6613 5485 6647
rect 5427 6607 5485 6613
rect 8460 6604 8466 6656
rect 8518 6644 8524 6656
rect 10116 6644 10122 6656
rect 8518 6616 10122 6644
rect 8518 6604 8524 6616
rect 10116 6604 10122 6616
rect 10174 6604 10180 6656
rect 1086 6554 58862 6576
rect 1086 6502 4228 6554
rect 4280 6502 4292 6554
rect 4344 6502 4356 6554
rect 4408 6502 4420 6554
rect 4472 6502 34948 6554
rect 35000 6502 35012 6554
rect 35064 6502 35076 6554
rect 35128 6502 35140 6554
rect 35192 6502 58862 6554
rect 1086 6480 58862 6502
rect 8184 6400 8190 6452
rect 8242 6440 8248 6452
rect 8460 6440 8466 6452
rect 8242 6400 8276 6440
rect 8248 6324 8276 6400
rect 8432 6400 8466 6440
rect 8518 6400 8524 6452
rect 17292 6440 17298 6452
rect 8616 6412 17298 6440
rect 8432 6324 8460 6400
rect 8616 6324 8644 6412
rect 17292 6400 17298 6412
rect 17350 6400 17356 6452
rect 18948 6304 18954 6316
rect 8814 6276 18954 6304
rect 18948 6264 18954 6276
rect 19006 6264 19012 6316
rect 10395 6239 10453 6245
rect 10395 6205 10407 6239
rect 10441 6205 10453 6239
rect 10395 6199 10453 6205
rect 10410 6168 10438 6199
rect 10576 6196 10582 6248
rect 10634 6236 10640 6248
rect 36523 6239 36581 6245
rect 36523 6236 36535 6239
rect 10634 6208 36535 6236
rect 10634 6196 10640 6208
rect 36523 6205 36535 6208
rect 36569 6205 36581 6239
rect 36523 6199 36581 6205
rect 26216 6168 26222 6180
rect 10410 6140 26222 6168
rect 26216 6128 26222 6140
rect 26274 6128 26280 6180
rect 14440 6100 14446 6112
rect 8906 6072 14446 6100
rect 14440 6060 14446 6072
rect 14498 6060 14504 6112
rect 1086 6010 58862 6032
rect 1086 5958 19588 6010
rect 19640 5958 19652 6010
rect 19704 5958 19716 6010
rect 19768 5958 19780 6010
rect 19832 5958 50308 6010
rect 50360 5958 50372 6010
rect 50424 5958 50436 6010
rect 50488 5958 50500 6010
rect 50552 5958 58862 6010
rect 1086 5936 58862 5958
rect 1284 5856 1290 5908
rect 1342 5896 1348 5908
rect 8460 5896 8466 5908
rect 1342 5868 8466 5896
rect 1342 5856 1348 5868
rect 8460 5856 8466 5868
rect 8518 5856 8524 5908
rect 20604 5856 20610 5908
rect 20662 5896 20668 5908
rect 28335 5899 28393 5905
rect 28335 5896 28347 5899
rect 20662 5868 28347 5896
rect 20662 5856 20668 5868
rect 28335 5865 28347 5868
rect 28381 5865 28393 5899
rect 28335 5859 28393 5865
rect 4596 5584 4602 5636
rect 4654 5624 4660 5636
rect 43515 5627 43573 5633
rect 43515 5624 43527 5627
rect 4654 5596 43527 5624
rect 4654 5584 4660 5596
rect 43515 5593 43527 5596
rect 43561 5593 43573 5627
rect 43515 5587 43573 5593
rect 14900 5516 14906 5568
rect 14958 5556 14964 5568
rect 18951 5559 19009 5565
rect 18951 5556 18963 5559
rect 14958 5528 18963 5556
rect 14958 5516 14964 5528
rect 18951 5525 18963 5528
rect 18997 5525 19009 5559
rect 18951 5519 19009 5525
rect 1086 5466 58862 5488
rect 1086 5414 4228 5466
rect 4280 5414 4292 5466
rect 4344 5414 4356 5466
rect 4408 5414 4420 5466
rect 4472 5414 34948 5466
rect 35000 5414 35012 5466
rect 35064 5414 35076 5466
rect 35128 5414 35140 5466
rect 35192 5414 58862 5466
rect 1086 5392 58862 5414
rect 12416 5352 12422 5364
rect 8432 5324 12422 5352
rect 8230 5210 8236 5262
rect 8288 5210 8294 5262
rect 8432 5236 8460 5324
rect 12416 5312 12422 5324
rect 12474 5312 12480 5364
rect 11312 5216 11318 5228
rect 8630 5188 11318 5216
rect 11312 5176 11318 5188
rect 11370 5176 11376 5228
rect 8736 5108 8742 5160
rect 8794 5148 8800 5160
rect 15268 5148 15274 5160
rect 8794 5120 15274 5148
rect 8794 5108 8800 5120
rect 15268 5108 15274 5120
rect 15326 5108 15332 5160
rect 8644 4972 8650 5024
rect 8702 4972 8708 5024
rect 20972 4972 20978 5024
rect 21030 5012 21036 5024
rect 21708 5012 21714 5024
rect 21030 4984 21714 5012
rect 21030 4972 21036 4984
rect 21708 4972 21714 4984
rect 21766 4972 21772 5024
rect 1086 4922 58862 4944
rect 1086 4870 19588 4922
rect 19640 4870 19652 4922
rect 19704 4870 19716 4922
rect 19768 4870 19780 4922
rect 19832 4870 50308 4922
rect 50360 4870 50372 4922
rect 50424 4870 50436 4922
rect 50488 4870 50500 4922
rect 50552 4870 58862 4922
rect 1086 4848 58862 4870
rect 12784 4768 12790 4820
rect 12842 4808 12848 4820
rect 12968 4808 12974 4820
rect 12842 4780 12974 4808
rect 12842 4768 12848 4780
rect 12968 4768 12974 4780
rect 13026 4768 13032 4820
rect 17016 4768 17022 4820
rect 17074 4808 17080 4820
rect 17384 4808 17390 4820
rect 17074 4780 17390 4808
rect 17074 4768 17080 4780
rect 17384 4768 17390 4780
rect 17442 4768 17448 4820
rect 40200 4768 40206 4820
rect 40258 4808 40264 4820
rect 41120 4808 41126 4820
rect 40258 4780 41126 4808
rect 40258 4768 40264 4780
rect 41120 4768 41126 4780
rect 41178 4768 41184 4820
rect 30080 4632 30086 4684
rect 30138 4672 30144 4684
rect 37256 4672 37262 4684
rect 30138 4644 37262 4672
rect 30138 4632 30144 4644
rect 37256 4632 37262 4644
rect 37314 4632 37320 4684
rect 23824 4496 23830 4548
rect 23882 4536 23888 4548
rect 31644 4536 31650 4548
rect 23882 4508 31650 4536
rect 23882 4496 23888 4508
rect 31644 4496 31650 4508
rect 31702 4496 31708 4548
rect 38268 4496 38274 4548
rect 38326 4536 38332 4548
rect 47008 4536 47014 4548
rect 38326 4508 47014 4536
rect 38326 4496 38332 4508
rect 47008 4496 47014 4508
rect 47066 4496 47072 4548
rect 7448 4428 7454 4480
rect 7506 4468 7512 4480
rect 31828 4468 31834 4480
rect 7506 4440 31834 4468
rect 7506 4428 7512 4440
rect 31828 4428 31834 4440
rect 31886 4428 31892 4480
rect 41028 4428 41034 4480
rect 41086 4468 41092 4480
rect 47655 4471 47713 4477
rect 47655 4468 47667 4471
rect 41086 4440 47667 4468
rect 41086 4428 41092 4440
rect 47655 4437 47667 4440
rect 47701 4437 47713 4471
rect 47655 4431 47713 4437
rect 1086 4378 58862 4400
rect 1086 4326 4228 4378
rect 4280 4326 4292 4378
rect 4344 4326 4356 4378
rect 4408 4326 4420 4378
rect 4472 4326 34948 4378
rect 35000 4326 35012 4378
rect 35064 4326 35076 4378
rect 35128 4326 35140 4378
rect 35192 4326 58862 4378
rect 1086 4304 58862 4326
rect 7448 4264 7454 4276
rect 7409 4236 7454 4264
rect 7448 4224 7454 4236
rect 7506 4224 7512 4276
rect 9104 4264 9110 4276
rect 8722 4236 9110 4264
rect 9104 4224 9110 4236
rect 9162 4224 9168 4276
rect 21156 4224 21162 4276
rect 21214 4264 21220 4276
rect 22260 4264 22266 4276
rect 21214 4236 22266 4264
rect 21214 4224 21220 4236
rect 22260 4224 22266 4236
rect 22318 4224 22324 4276
rect 25020 4224 25026 4276
rect 25078 4264 25084 4276
rect 43144 4264 43150 4276
rect 25078 4236 29758 4264
rect 25078 4224 25084 4236
rect 18948 4156 18954 4208
rect 19006 4196 19012 4208
rect 27412 4196 27418 4208
rect 19006 4168 27418 4196
rect 19006 4156 19012 4168
rect 27412 4156 27418 4168
rect 27470 4156 27476 4208
rect 3676 4088 3682 4140
rect 3734 4128 3740 4140
rect 3952 4128 3958 4140
rect 3734 4100 3958 4128
rect 3734 4088 3740 4100
rect 3952 4088 3958 4100
rect 4010 4088 4016 4140
rect 4688 4088 4694 4140
rect 4746 4128 4752 4140
rect 5148 4128 5154 4140
rect 4746 4100 5154 4128
rect 4746 4088 4752 4100
rect 5148 4088 5154 4100
rect 5206 4088 5212 4140
rect 6160 4088 6166 4140
rect 6218 4128 6224 4140
rect 6712 4128 6718 4140
rect 6218 4100 6718 4128
rect 6218 4088 6224 4100
rect 6712 4088 6718 4100
rect 6770 4088 6776 4140
rect 7632 4088 7638 4140
rect 7690 4128 7696 4140
rect 8000 4128 8006 4140
rect 7690 4100 8006 4128
rect 7690 4088 7696 4100
rect 8000 4088 8006 4100
rect 8058 4088 8064 4140
rect 8092 4088 8098 4140
rect 8150 4128 8156 4140
rect 8150 4100 8262 4128
rect 8150 4088 8156 4100
rect 9840 4088 9846 4140
rect 9898 4128 9904 4140
rect 10760 4128 10766 4140
rect 9898 4100 10766 4128
rect 9898 4088 9904 4100
rect 10760 4088 10766 4100
rect 10818 4088 10824 4140
rect 11680 4088 11686 4140
rect 11738 4128 11744 4140
rect 12324 4128 12330 4140
rect 11738 4100 12330 4128
rect 11738 4088 11744 4100
rect 12324 4088 12330 4100
rect 12382 4088 12388 4140
rect 13060 4088 13066 4140
rect 13118 4128 13124 4140
rect 13336 4128 13342 4140
rect 13118 4100 13342 4128
rect 13118 4088 13124 4100
rect 13336 4088 13342 4100
rect 13394 4088 13400 4140
rect 13428 4088 13434 4140
rect 13486 4128 13492 4140
rect 13704 4128 13710 4140
rect 13486 4100 13710 4128
rect 13486 4088 13492 4100
rect 13704 4088 13710 4100
rect 13762 4088 13768 4140
rect 14532 4088 14538 4140
rect 14590 4128 14596 4140
rect 15452 4128 15458 4140
rect 14590 4100 15458 4128
rect 14590 4088 14596 4100
rect 15452 4088 15458 4100
rect 15510 4088 15516 4140
rect 16004 4088 16010 4140
rect 16062 4128 16068 4140
rect 16464 4128 16470 4140
rect 16062 4100 16470 4128
rect 16062 4088 16068 4100
rect 16464 4088 16470 4100
rect 16522 4088 16528 4140
rect 17108 4088 17114 4140
rect 17166 4128 17172 4140
rect 17844 4128 17850 4140
rect 17166 4100 17850 4128
rect 17166 4088 17172 4100
rect 17844 4088 17850 4100
rect 17902 4088 17908 4140
rect 18856 4088 18862 4140
rect 18914 4128 18920 4140
rect 19316 4128 19322 4140
rect 18914 4100 19322 4128
rect 18914 4088 18920 4100
rect 19316 4088 19322 4100
rect 19374 4088 19380 4140
rect 20052 4088 20058 4140
rect 20110 4128 20116 4140
rect 20420 4128 20426 4140
rect 20110 4100 20426 4128
rect 20110 4088 20116 4100
rect 20420 4088 20426 4100
rect 20478 4088 20484 4140
rect 21248 4088 21254 4140
rect 21306 4128 21312 4140
rect 22628 4128 22634 4140
rect 21306 4100 22634 4128
rect 21306 4088 21312 4100
rect 22628 4088 22634 4100
rect 22686 4088 22692 4140
rect 24284 4088 24290 4140
rect 24342 4128 24348 4140
rect 25020 4128 25026 4140
rect 24342 4100 25026 4128
rect 24342 4088 24348 4100
rect 25020 4088 25026 4100
rect 25078 4088 25084 4140
rect 25204 4088 25210 4140
rect 25262 4128 25268 4140
rect 26124 4128 26130 4140
rect 25262 4100 26130 4128
rect 25262 4088 25268 4100
rect 26124 4088 26130 4100
rect 26182 4088 26188 4140
rect 26308 4088 26314 4140
rect 26366 4128 26372 4140
rect 27504 4128 27510 4140
rect 26366 4100 27510 4128
rect 26366 4088 26372 4100
rect 27504 4088 27510 4100
rect 27562 4088 27568 4140
rect 28516 4088 28522 4140
rect 28574 4128 28580 4140
rect 29620 4128 29626 4140
rect 28574 4100 29626 4128
rect 28574 4088 28580 4100
rect 29620 4088 29626 4100
rect 29678 4088 29684 4140
rect 29730 4128 29758 4236
rect 37734 4236 43150 4264
rect 30558 4168 31414 4196
rect 30558 4128 30586 4168
rect 29730 4100 30586 4128
rect 31386 4128 31414 4168
rect 31386 4100 31598 4128
rect 3216 4020 3222 4072
rect 3274 4060 3280 4072
rect 4044 4060 4050 4072
rect 3274 4032 4050 4060
rect 3274 4020 3280 4032
rect 4044 4020 4050 4032
rect 4102 4020 4108 4072
rect 5056 4020 5062 4072
rect 5114 4060 5120 4072
rect 5424 4060 5430 4072
rect 5114 4032 5430 4060
rect 5114 4020 5120 4032
rect 5424 4020 5430 4032
rect 5482 4020 5488 4072
rect 11312 4020 11318 4072
rect 11370 4060 11376 4072
rect 12048 4060 12054 4072
rect 11370 4032 12054 4060
rect 11370 4020 11376 4032
rect 12048 4020 12054 4032
rect 12106 4020 12112 4072
rect 13796 4020 13802 4072
rect 13854 4060 13860 4072
rect 14992 4060 14998 4072
rect 13854 4032 14998 4060
rect 13854 4020 13860 4032
rect 14992 4020 14998 4032
rect 15050 4020 15056 4072
rect 19960 4020 19966 4072
rect 20018 4060 20024 4072
rect 20788 4060 20794 4072
rect 20018 4032 20794 4060
rect 20018 4020 20024 4032
rect 20788 4020 20794 4032
rect 20846 4020 20852 4072
rect 22812 4020 22818 4072
rect 22870 4060 22876 4072
rect 24836 4060 24842 4072
rect 22870 4032 24842 4060
rect 22870 4020 22876 4032
rect 24836 4020 24842 4032
rect 24894 4020 24900 4072
rect 27044 4020 27050 4072
rect 27102 4060 27108 4072
rect 27102 4032 28286 4060
rect 27102 4020 27108 4032
rect 4964 3952 4970 4004
rect 5022 3992 5028 4004
rect 6896 3992 6902 4004
rect 5022 3964 6902 3992
rect 5022 3952 5028 3964
rect 6896 3952 6902 3964
rect 6954 3952 6960 4004
rect 6252 3884 6258 3936
rect 6310 3924 6316 3936
rect 8432 3924 8460 4012
rect 12784 3952 12790 4004
rect 12842 3992 12848 4004
rect 13520 3992 13526 4004
rect 12842 3964 13526 3992
rect 12842 3952 12848 3964
rect 13520 3952 13526 3964
rect 13578 3952 13584 4004
rect 16832 3952 16838 4004
rect 16890 3992 16896 4004
rect 17844 3992 17850 4004
rect 16890 3964 17850 3992
rect 16890 3952 16896 3964
rect 17844 3952 17850 3964
rect 17902 3952 17908 4004
rect 20144 3952 20150 4004
rect 20202 3992 20208 4004
rect 21156 3992 21162 4004
rect 20202 3964 21162 3992
rect 20202 3952 20208 3964
rect 21156 3952 21162 3964
rect 21214 3952 21220 4004
rect 21248 3952 21254 4004
rect 21306 3992 21312 4004
rect 22536 3992 22542 4004
rect 21306 3964 22542 3992
rect 21306 3952 21312 3964
rect 22536 3952 22542 3964
rect 22594 3952 22600 4004
rect 25480 3952 25486 4004
rect 25538 3992 25544 4004
rect 28148 3992 28154 4004
rect 25538 3964 28154 3992
rect 25538 3952 25544 3964
rect 28148 3952 28154 3964
rect 28206 3952 28212 4004
rect 28258 3992 28286 4032
rect 28884 4020 28890 4072
rect 28942 4060 28948 4072
rect 30172 4060 30178 4072
rect 28942 4032 30178 4060
rect 28942 4020 28948 4032
rect 30172 4020 30178 4032
rect 30230 4020 30236 4072
rect 31570 4060 31598 4100
rect 31644 4088 31650 4140
rect 31702 4128 31708 4140
rect 37734 4128 37762 4236
rect 43144 4224 43150 4236
rect 43202 4224 43208 4276
rect 31702 4100 37762 4128
rect 37826 4168 38774 4196
rect 31702 4088 31708 4100
rect 31570 4032 33898 4060
rect 32840 3992 32846 4004
rect 28258 3964 32846 3992
rect 32840 3952 32846 3964
rect 32898 3952 32904 4004
rect 33870 3992 33898 4032
rect 33944 4020 33950 4072
rect 34002 4060 34008 4072
rect 34404 4060 34410 4072
rect 34002 4032 34410 4060
rect 34002 4020 34008 4032
rect 34404 4020 34410 4032
rect 34462 4020 34468 4072
rect 34588 4020 34594 4072
rect 34646 4060 34652 4072
rect 37826 4060 37854 4168
rect 34646 4032 37854 4060
rect 34646 4020 34652 4032
rect 37992 4020 37998 4072
rect 38050 4060 38056 4072
rect 38544 4060 38550 4072
rect 38050 4032 38550 4060
rect 38050 4020 38056 4032
rect 38544 4020 38550 4032
rect 38602 4020 38608 4072
rect 38746 4060 38774 4168
rect 39648 4156 39654 4208
rect 39706 4196 39712 4208
rect 39706 4168 46870 4196
rect 39706 4156 39712 4168
rect 46732 4128 46738 4140
rect 41598 4100 46738 4128
rect 39740 4060 39746 4072
rect 38746 4032 39746 4060
rect 39740 4020 39746 4032
rect 39798 4020 39804 4072
rect 41598 4060 41626 4100
rect 46732 4088 46738 4100
rect 46790 4088 46796 4140
rect 46842 4128 46870 4168
rect 50780 4128 50786 4140
rect 46842 4100 50786 4128
rect 50780 4088 50786 4100
rect 50838 4088 50844 4140
rect 51792 4088 51798 4140
rect 51850 4128 51856 4140
rect 54184 4128 54190 4140
rect 51850 4100 54190 4128
rect 51850 4088 51856 4100
rect 54184 4088 54190 4100
rect 54242 4088 54248 4140
rect 51608 4060 51614 4072
rect 41230 4032 41626 4060
rect 46198 4032 51614 4060
rect 41230 3992 41258 4032
rect 33870 3964 41258 3992
rect 6310 3896 8460 3924
rect 6310 3884 6316 3896
rect 10668 3884 10674 3936
rect 10726 3924 10732 3936
rect 14440 3924 14446 3936
rect 10726 3896 14446 3924
rect 10726 3884 10732 3896
rect 14440 3884 14446 3896
rect 14498 3884 14504 3936
rect 15728 3884 15734 3936
rect 15786 3924 15792 3936
rect 31736 3924 31742 3936
rect 15786 3896 31742 3924
rect 15786 3884 15792 3896
rect 31736 3884 31742 3896
rect 31794 3884 31800 3936
rect 31828 3884 31834 3936
rect 31886 3924 31892 3936
rect 33208 3924 33214 3936
rect 31886 3896 33214 3924
rect 31886 3884 31892 3896
rect 33208 3884 33214 3896
rect 33266 3884 33272 3936
rect 35232 3884 35238 3936
rect 35290 3924 35296 3936
rect 36520 3924 36526 3936
rect 35290 3896 36526 3924
rect 35290 3884 35296 3896
rect 36520 3884 36526 3896
rect 36578 3884 36584 3936
rect 36612 3884 36618 3936
rect 36670 3924 36676 3936
rect 39096 3924 39102 3936
rect 36670 3896 39102 3924
rect 36670 3884 36676 3896
rect 39096 3884 39102 3896
rect 39154 3884 39160 3936
rect 39188 3884 39194 3936
rect 39246 3924 39252 3936
rect 40568 3924 40574 3936
rect 39246 3896 40574 3924
rect 39246 3884 39252 3896
rect 40568 3884 40574 3896
rect 40626 3884 40632 3936
rect 40752 3884 40758 3936
rect 40810 3924 40816 3936
rect 46198 3924 46226 4032
rect 51608 4020 51614 4032
rect 51666 4020 51672 4072
rect 49768 3952 49774 4004
rect 49826 3992 49832 4004
rect 50964 3992 50970 4004
rect 49826 3964 50970 3992
rect 49826 3952 49832 3964
rect 50964 3952 50970 3964
rect 51022 3952 51028 4004
rect 40810 3896 46226 3924
rect 40810 3884 40816 3896
rect 48940 3884 48946 3936
rect 48998 3924 49004 3936
rect 56760 3924 56766 3936
rect 48998 3896 56766 3924
rect 48998 3884 49004 3896
rect 56760 3884 56766 3896
rect 56818 3884 56824 3936
rect 1086 3834 58862 3856
rect 1086 3782 19588 3834
rect 19640 3782 19652 3834
rect 19704 3782 19716 3834
rect 19768 3782 19780 3834
rect 19832 3782 50308 3834
rect 50360 3782 50372 3834
rect 50424 3782 50436 3834
rect 50488 3782 50500 3834
rect 50552 3782 58862 3834
rect 1086 3760 58862 3782
rect 8368 3680 8374 3732
rect 8426 3720 8432 3732
rect 11772 3720 11778 3732
rect 8426 3692 11778 3720
rect 8426 3680 8432 3692
rect 11772 3680 11778 3692
rect 11830 3680 11836 3732
rect 11864 3680 11870 3732
rect 11922 3720 11928 3732
rect 11922 3692 19178 3720
rect 11922 3680 11928 3692
rect 7264 3612 7270 3664
rect 7322 3652 7328 3664
rect 11036 3652 11042 3664
rect 7322 3624 11042 3652
rect 7322 3612 7328 3624
rect 11036 3612 11042 3624
rect 11094 3612 11100 3664
rect 12876 3612 12882 3664
rect 12934 3652 12940 3664
rect 14808 3652 14814 3664
rect 12934 3624 14814 3652
rect 12934 3612 12940 3624
rect 14808 3612 14814 3624
rect 14866 3612 14872 3664
rect 19150 3652 19178 3692
rect 23180 3680 23186 3732
rect 23238 3720 23244 3732
rect 24284 3720 24290 3732
rect 23238 3692 24290 3720
rect 23238 3680 23244 3692
rect 24284 3680 24290 3692
rect 24342 3680 24348 3732
rect 27504 3680 27510 3732
rect 27562 3720 27568 3732
rect 28976 3720 28982 3732
rect 27562 3692 28982 3720
rect 27562 3680 27568 3692
rect 28976 3680 28982 3692
rect 29034 3680 29040 3732
rect 31736 3680 31742 3732
rect 31794 3720 31800 3732
rect 32932 3720 32938 3732
rect 31794 3692 32938 3720
rect 31794 3680 31800 3692
rect 32932 3680 32938 3692
rect 32990 3680 32996 3732
rect 33024 3680 33030 3732
rect 33082 3720 33088 3732
rect 39188 3720 39194 3732
rect 33082 3692 39194 3720
rect 33082 3680 33088 3692
rect 39188 3680 39194 3692
rect 39246 3680 39252 3732
rect 48664 3720 48670 3732
rect 41598 3692 48670 3720
rect 31828 3652 31834 3664
rect 19150 3624 31834 3652
rect 31828 3612 31834 3624
rect 31886 3612 31892 3664
rect 40384 3652 40390 3664
rect 36538 3624 40390 3652
rect 180 3544 186 3596
rect 238 3584 244 3596
rect 1008 3584 1014 3596
rect 238 3556 1014 3584
rect 238 3544 244 3556
rect 1008 3544 1014 3556
rect 1066 3544 1072 3596
rect 1376 3544 1382 3596
rect 1434 3584 1440 3596
rect 2388 3584 2394 3596
rect 1434 3556 2394 3584
rect 1434 3544 1440 3556
rect 2388 3544 2394 3556
rect 2446 3544 2452 3596
rect 6344 3544 6350 3596
rect 6402 3584 6408 3596
rect 14348 3584 14354 3596
rect 6402 3556 14354 3584
rect 6402 3544 6408 3556
rect 14348 3544 14354 3556
rect 14406 3544 14412 3596
rect 17292 3544 17298 3596
rect 17350 3584 17356 3596
rect 36538 3584 36566 3624
rect 40384 3612 40390 3624
rect 40442 3612 40448 3664
rect 17350 3556 36566 3584
rect 17350 3544 17356 3556
rect 36612 3544 36618 3596
rect 36670 3584 36676 3596
rect 38636 3584 38642 3596
rect 36670 3556 38642 3584
rect 36670 3544 36676 3556
rect 38636 3544 38642 3556
rect 38694 3544 38700 3596
rect 38728 3544 38734 3596
rect 38786 3584 38792 3596
rect 39924 3584 39930 3596
rect 38786 3556 39930 3584
rect 38786 3544 38792 3556
rect 39924 3544 39930 3556
rect 39982 3544 39988 3596
rect 5332 3476 5338 3528
rect 5390 3516 5396 3528
rect 31644 3516 31650 3528
rect 5390 3488 31650 3516
rect 5390 3476 5396 3488
rect 31644 3476 31650 3488
rect 31702 3476 31708 3528
rect 31754 3488 31966 3516
rect 3032 3408 3038 3460
rect 3090 3448 3096 3460
rect 31754 3448 31782 3488
rect 3090 3420 31782 3448
rect 31938 3448 31966 3488
rect 37808 3476 37814 3528
rect 37866 3516 37872 3528
rect 41598 3516 41626 3692
rect 48664 3680 48670 3692
rect 48722 3680 48728 3732
rect 49032 3680 49038 3732
rect 49090 3720 49096 3732
rect 49090 3692 51654 3720
rect 49090 3680 49096 3692
rect 42040 3612 42046 3664
rect 42098 3652 42104 3664
rect 46916 3652 46922 3664
rect 42098 3624 46922 3652
rect 42098 3612 42104 3624
rect 46916 3612 46922 3624
rect 46974 3612 46980 3664
rect 47468 3612 47474 3664
rect 47526 3652 47532 3664
rect 49952 3652 49958 3664
rect 47526 3624 49958 3652
rect 47526 3612 47532 3624
rect 49952 3612 49958 3624
rect 50010 3612 50016 3664
rect 51240 3652 51246 3664
rect 50062 3624 51246 3652
rect 47928 3544 47934 3596
rect 47986 3584 47992 3596
rect 50062 3584 50090 3624
rect 51240 3612 51246 3624
rect 51298 3612 51304 3664
rect 51626 3652 51654 3692
rect 51700 3680 51706 3732
rect 51758 3720 51764 3732
rect 59336 3720 59342 3732
rect 51758 3692 59342 3720
rect 51758 3680 51764 3692
rect 59336 3680 59342 3692
rect 59394 3680 59400 3732
rect 57496 3652 57502 3664
rect 51626 3624 57502 3652
rect 57496 3612 57502 3624
rect 57554 3612 57560 3664
rect 47986 3556 50090 3584
rect 47986 3544 47992 3556
rect 50136 3544 50142 3596
rect 50194 3584 50200 3596
rect 54920 3584 54926 3596
rect 50194 3556 54926 3584
rect 50194 3544 50200 3556
rect 54920 3544 54926 3556
rect 54978 3544 54984 3596
rect 37866 3488 41626 3516
rect 37866 3476 37872 3488
rect 47284 3476 47290 3528
rect 47342 3516 47348 3528
rect 48296 3516 48302 3528
rect 47342 3488 48302 3516
rect 47342 3476 47348 3488
rect 48296 3476 48302 3488
rect 48354 3476 48360 3528
rect 53816 3516 53822 3528
rect 50890 3488 53822 3516
rect 39924 3448 39930 3460
rect 31938 3420 39930 3448
rect 3090 3408 3096 3420
rect 39924 3408 39930 3420
rect 39982 3408 39988 3460
rect 45720 3408 45726 3460
rect 45778 3448 45784 3460
rect 46824 3448 46830 3460
rect 45778 3420 46830 3448
rect 45778 3408 45784 3420
rect 46824 3408 46830 3420
rect 46882 3408 46888 3460
rect 47008 3408 47014 3460
rect 47066 3448 47072 3460
rect 50890 3448 50918 3488
rect 53816 3476 53822 3488
rect 53874 3476 53880 3528
rect 47066 3420 50918 3448
rect 47066 3408 47072 3420
rect 14624 3340 14630 3392
rect 14682 3380 14688 3392
rect 21248 3380 21254 3392
rect 14682 3352 21254 3380
rect 14682 3340 14688 3352
rect 21248 3340 21254 3352
rect 21306 3340 21312 3392
rect 21432 3340 21438 3392
rect 21490 3380 21496 3392
rect 22076 3380 22082 3392
rect 21490 3352 22082 3380
rect 21490 3340 21496 3352
rect 22076 3340 22082 3352
rect 22134 3340 22140 3392
rect 23088 3340 23094 3392
rect 23146 3380 23152 3392
rect 23916 3380 23922 3392
rect 23146 3352 23922 3380
rect 23146 3340 23152 3352
rect 23916 3340 23922 3352
rect 23974 3340 23980 3392
rect 24376 3340 24382 3392
rect 24434 3380 24440 3392
rect 27044 3380 27050 3392
rect 24434 3352 27050 3380
rect 24434 3340 24440 3352
rect 27044 3340 27050 3352
rect 27102 3340 27108 3392
rect 28332 3340 28338 3392
rect 28390 3380 28396 3392
rect 31092 3380 31098 3392
rect 28390 3352 31098 3380
rect 28390 3340 28396 3352
rect 31092 3340 31098 3352
rect 31150 3340 31156 3392
rect 31644 3340 31650 3392
rect 31702 3380 31708 3392
rect 34588 3380 34594 3392
rect 31702 3352 34594 3380
rect 31702 3340 31708 3352
rect 34588 3340 34594 3352
rect 34646 3340 34652 3392
rect 36520 3340 36526 3392
rect 36578 3380 36584 3392
rect 46088 3380 46094 3392
rect 36578 3352 46094 3380
rect 36578 3340 36584 3352
rect 46088 3340 46094 3352
rect 46146 3340 46152 3392
rect 47560 3340 47566 3392
rect 47618 3380 47624 3392
rect 52347 3383 52405 3389
rect 52347 3380 52359 3383
rect 47618 3352 52359 3380
rect 47618 3340 47624 3352
rect 52347 3349 52359 3352
rect 52393 3349 52405 3383
rect 52347 3343 52405 3349
rect 55288 3340 55294 3392
rect 55346 3380 55352 3392
rect 58419 3383 58477 3389
rect 58419 3380 58431 3383
rect 55346 3352 58431 3380
rect 55346 3340 55352 3352
rect 58419 3349 58431 3352
rect 58465 3349 58477 3383
rect 58419 3343 58477 3349
rect 1086 3290 58862 3312
rect 1086 3238 4228 3290
rect 4280 3238 4292 3290
rect 4344 3238 4356 3290
rect 4408 3238 4420 3290
rect 4472 3238 34948 3290
rect 35000 3238 35012 3290
rect 35064 3238 35076 3290
rect 35128 3238 35140 3290
rect 35192 3238 58862 3290
rect 1086 3216 58862 3238
rect 6068 3136 6074 3188
rect 6126 3176 6132 3188
rect 6126 3148 8722 3176
rect 6126 3136 6132 3148
rect 10852 3136 10858 3188
rect 10910 3176 10916 3188
rect 17292 3176 17298 3188
rect 10910 3148 17298 3176
rect 10910 3136 10916 3148
rect 17292 3136 17298 3148
rect 17350 3136 17356 3188
rect 18580 3176 18586 3188
rect 18541 3148 18586 3176
rect 18580 3136 18586 3148
rect 18638 3136 18644 3188
rect 22536 3136 22542 3188
rect 22594 3176 22600 3188
rect 36152 3176 36158 3188
rect 22594 3148 36158 3176
rect 22594 3136 22600 3148
rect 36152 3136 36158 3148
rect 36210 3136 36216 3188
rect 38360 3136 38366 3188
rect 38418 3176 38424 3188
rect 41028 3176 41034 3188
rect 38418 3148 41034 3176
rect 38418 3136 38424 3148
rect 41028 3136 41034 3148
rect 41086 3136 41092 3188
rect 41304 3136 41310 3188
rect 41362 3176 41368 3188
rect 45260 3176 45266 3188
rect 41362 3148 45266 3176
rect 41362 3136 41368 3148
rect 45260 3136 45266 3148
rect 45318 3136 45324 3188
rect 46916 3136 46922 3188
rect 46974 3176 46980 3188
rect 50136 3176 50142 3188
rect 46974 3148 50142 3176
rect 46974 3136 46980 3148
rect 50136 3136 50142 3148
rect 50194 3136 50200 3188
rect 50596 3136 50602 3188
rect 50654 3176 50660 3188
rect 58968 3176 58974 3188
rect 50654 3148 58974 3176
rect 50654 3136 50660 3148
rect 58968 3136 58974 3148
rect 59026 3136 59032 3188
rect 8828 3068 8834 3120
rect 8886 3108 8892 3120
rect 19040 3108 19046 3120
rect 8886 3080 19046 3108
rect 8886 3068 8892 3080
rect 19040 3068 19046 3080
rect 19098 3068 19104 3120
rect 23364 3068 23370 3120
rect 23422 3108 23428 3120
rect 25940 3108 25946 3120
rect 23422 3080 25946 3108
rect 23422 3068 23428 3080
rect 25940 3068 25946 3080
rect 25998 3068 26004 3120
rect 26952 3068 26958 3120
rect 27010 3108 27016 3120
rect 29620 3108 29626 3120
rect 27010 3080 29626 3108
rect 27010 3068 27016 3080
rect 29620 3068 29626 3080
rect 29678 3068 29684 3120
rect 38084 3068 38090 3120
rect 38142 3108 38148 3120
rect 47928 3108 47934 3120
rect 38142 3080 47934 3108
rect 38142 3068 38148 3080
rect 47928 3068 47934 3080
rect 47986 3068 47992 3120
rect 49676 3068 49682 3120
rect 49734 3108 49740 3120
rect 50504 3108 50510 3120
rect 49734 3080 50510 3108
rect 49734 3068 49740 3080
rect 50504 3068 50510 3080
rect 50562 3068 50568 3120
rect 50688 3068 50694 3120
rect 50746 3108 50752 3120
rect 58232 3108 58238 3120
rect 50746 3080 58238 3108
rect 50746 3068 50752 3080
rect 58232 3068 58238 3080
rect 58290 3068 58296 3120
rect 2664 3000 2670 3052
rect 2722 3040 2728 3052
rect 2722 3012 8262 3040
rect 2722 3000 2728 3012
rect 8460 3000 8466 3052
rect 8518 3000 8524 3052
rect 16280 3000 16286 3052
rect 16338 3040 16344 3052
rect 18580 3040 18586 3052
rect 16338 3012 18586 3040
rect 16338 3000 16344 3012
rect 18580 3000 18586 3012
rect 18638 3000 18644 3052
rect 21064 3000 21070 3052
rect 21122 3040 21128 3052
rect 23732 3040 23738 3052
rect 21122 3012 23738 3040
rect 21122 3000 21128 3012
rect 23732 3000 23738 3012
rect 23790 3000 23796 3052
rect 24192 3000 24198 3052
rect 24250 3040 24256 3052
rect 27412 3040 27418 3052
rect 24250 3012 27418 3040
rect 24250 3000 24256 3012
rect 27412 3000 27418 3012
rect 27470 3000 27476 3052
rect 27872 3000 27878 3052
rect 27930 3040 27936 3052
rect 28332 3040 28338 3052
rect 27930 3012 28338 3040
rect 27930 3000 27936 3012
rect 28332 3000 28338 3012
rect 28390 3000 28396 3052
rect 29528 3000 29534 3052
rect 29586 3040 29592 3052
rect 36520 3040 36526 3052
rect 29586 3012 36526 3040
rect 29586 3000 29592 3012
rect 36520 3000 36526 3012
rect 36578 3000 36584 3052
rect 38176 3000 38182 3052
rect 38234 3040 38240 3052
rect 38234 3012 39602 3040
rect 38234 3000 38240 3012
rect 8478 2972 8506 3000
rect 8446 2944 8506 2972
rect 20696 2932 20702 2984
rect 20754 2972 20760 2984
rect 23364 2972 23370 2984
rect 20754 2944 23370 2972
rect 20754 2932 20760 2944
rect 23364 2932 23370 2944
rect 23422 2932 23428 2984
rect 26216 2932 26222 2984
rect 26274 2972 26280 2984
rect 29344 2972 29350 2984
rect 26274 2944 29350 2972
rect 26274 2932 26280 2944
rect 29344 2932 29350 2944
rect 29402 2932 29408 2984
rect 29436 2932 29442 2984
rect 29494 2972 29500 2984
rect 39464 2972 39470 2984
rect 29494 2944 39470 2972
rect 29494 2932 29500 2944
rect 39464 2932 39470 2944
rect 39522 2932 39528 2984
rect 39574 2972 39602 3012
rect 39740 3000 39746 3052
rect 39798 3040 39804 3052
rect 41212 3040 41218 3052
rect 39798 3012 41218 3040
rect 39798 3000 39804 3012
rect 41212 3000 41218 3012
rect 41270 3000 41276 3052
rect 41396 3000 41402 3052
rect 41454 3040 41460 3052
rect 51976 3040 51982 3052
rect 41454 3012 51982 3040
rect 41454 3000 41460 3012
rect 51976 3000 51982 3012
rect 52034 3000 52040 3052
rect 54552 3000 54558 3052
rect 54610 3040 54616 3052
rect 55104 3040 55110 3052
rect 54610 3012 55110 3040
rect 54610 3000 54616 3012
rect 55104 3000 55110 3012
rect 55162 3000 55168 3052
rect 42776 2972 42782 2984
rect 39574 2944 42782 2972
rect 42776 2932 42782 2944
rect 42834 2932 42840 2984
rect 45260 2932 45266 2984
rect 45318 2972 45324 2984
rect 49032 2972 49038 2984
rect 45318 2944 49038 2972
rect 45318 2932 45324 2944
rect 49032 2932 49038 2944
rect 49090 2932 49096 2984
rect 56392 2972 56398 2984
rect 49142 2944 56398 2972
rect 22352 2864 22358 2916
rect 22410 2904 22416 2916
rect 26676 2904 26682 2916
rect 22410 2876 26682 2904
rect 22410 2864 22416 2876
rect 26676 2864 26682 2876
rect 26734 2864 26740 2916
rect 28424 2864 28430 2916
rect 28482 2904 28488 2916
rect 28482 2876 30954 2904
rect 28482 2864 28488 2876
rect 9564 2796 9570 2848
rect 9622 2836 9628 2848
rect 12048 2836 12054 2848
rect 9622 2808 12054 2836
rect 9622 2796 9628 2808
rect 12048 2796 12054 2808
rect 12106 2796 12112 2848
rect 27136 2796 27142 2848
rect 27194 2836 27200 2848
rect 30816 2836 30822 2848
rect 27194 2808 30822 2836
rect 27194 2796 27200 2808
rect 30816 2796 30822 2808
rect 30874 2796 30880 2848
rect 30926 2836 30954 2876
rect 31092 2864 31098 2916
rect 31150 2904 31156 2916
rect 33576 2904 33582 2916
rect 31150 2876 33582 2904
rect 31150 2864 31156 2876
rect 33576 2864 33582 2876
rect 33634 2864 33640 2916
rect 33668 2864 33674 2916
rect 33726 2904 33732 2916
rect 33726 2876 34450 2904
rect 33726 2864 33732 2876
rect 34312 2836 34318 2848
rect 30926 2808 34318 2836
rect 34312 2796 34318 2808
rect 34370 2796 34376 2848
rect 34422 2836 34450 2876
rect 34588 2864 34594 2916
rect 34646 2904 34652 2916
rect 39832 2904 39838 2916
rect 34646 2876 39838 2904
rect 34646 2864 34652 2876
rect 39832 2864 39838 2876
rect 39890 2864 39896 2916
rect 41304 2864 41310 2916
rect 41362 2904 41368 2916
rect 41672 2904 41678 2916
rect 41362 2876 41678 2904
rect 41362 2864 41368 2876
rect 41672 2864 41678 2876
rect 41730 2864 41736 2916
rect 42132 2864 42138 2916
rect 42190 2904 42196 2916
rect 42190 2876 44386 2904
rect 42190 2864 42196 2876
rect 40752 2836 40758 2848
rect 34422 2808 40758 2836
rect 40752 2796 40758 2808
rect 40810 2796 40816 2848
rect 40844 2796 40850 2848
rect 40902 2836 40908 2848
rect 44248 2836 44254 2848
rect 40902 2808 44254 2836
rect 40902 2796 40908 2808
rect 44248 2796 44254 2808
rect 44306 2796 44312 2848
rect 44358 2836 44386 2876
rect 44800 2864 44806 2916
rect 44858 2904 44864 2916
rect 49142 2904 49170 2944
rect 56392 2932 56398 2944
rect 56450 2932 56456 2984
rect 44858 2876 49170 2904
rect 44858 2864 44864 2876
rect 50780 2864 50786 2916
rect 50838 2904 50844 2916
rect 53448 2904 53454 2916
rect 50838 2876 53454 2904
rect 50838 2864 50844 2876
rect 53448 2864 53454 2876
rect 53506 2864 53512 2916
rect 49676 2836 49682 2848
rect 44358 2808 49682 2836
rect 49676 2796 49682 2808
rect 49734 2796 49740 2848
rect 50044 2796 50050 2848
rect 50102 2836 50108 2848
rect 57864 2836 57870 2848
rect 50102 2808 57870 2836
rect 50102 2796 50108 2808
rect 57864 2796 57870 2808
rect 57922 2796 57928 2848
rect 1086 2746 58862 2768
rect 1086 2694 19588 2746
rect 19640 2694 19652 2746
rect 19704 2694 19716 2746
rect 19768 2694 19780 2746
rect 19832 2694 50308 2746
rect 50360 2694 50372 2746
rect 50424 2694 50436 2746
rect 50488 2694 50500 2746
rect 50552 2694 58862 2746
rect 1086 2672 58862 2694
rect 22444 2592 22450 2644
rect 22502 2632 22508 2644
rect 22812 2632 22818 2644
rect 22502 2604 22818 2632
rect 22502 2592 22508 2604
rect 22812 2592 22818 2604
rect 22870 2592 22876 2644
rect 22904 2592 22910 2644
rect 22962 2632 22968 2644
rect 23180 2632 23186 2644
rect 22962 2604 23186 2632
rect 22962 2592 22968 2604
rect 23180 2592 23186 2604
rect 23238 2592 23244 2644
rect 25664 2592 25670 2644
rect 25722 2632 25728 2644
rect 27780 2632 27786 2644
rect 25722 2604 27786 2632
rect 25722 2592 25728 2604
rect 27780 2592 27786 2604
rect 27838 2592 27844 2644
rect 30816 2592 30822 2644
rect 30874 2632 30880 2644
rect 32472 2632 32478 2644
rect 30874 2604 32478 2632
rect 30874 2592 30880 2604
rect 32472 2592 32478 2604
rect 32530 2592 32536 2644
rect 39924 2592 39930 2644
rect 39982 2632 39988 2644
rect 40844 2632 40850 2644
rect 39982 2604 40850 2632
rect 39982 2592 39988 2604
rect 40844 2592 40850 2604
rect 40902 2592 40908 2644
rect 40384 2524 40390 2576
rect 40442 2564 40448 2576
rect 42408 2564 42414 2576
rect 40442 2536 42414 2564
rect 40442 2524 40448 2536
rect 42408 2524 42414 2536
rect 42466 2524 42472 2576
rect 48480 2524 48486 2576
rect 48538 2564 48544 2576
rect 53080 2564 53086 2576
rect 48538 2536 53086 2564
rect 48538 2524 48544 2536
rect 53080 2524 53086 2536
rect 53138 2524 53144 2576
rect 7359 2499 7417 2505
rect 7359 2465 7371 2499
rect 7405 2496 7417 2499
rect 9564 2496 9570 2508
rect 7405 2468 9570 2496
rect 7405 2465 7417 2468
rect 7359 2459 7417 2465
rect 9564 2456 9570 2468
rect 9622 2456 9628 2508
rect 12416 2456 12422 2508
rect 12474 2496 12480 2508
rect 13152 2496 13158 2508
rect 12474 2468 13158 2496
rect 12474 2456 12480 2468
rect 13152 2456 13158 2468
rect 13210 2456 13216 2508
rect 19411 2363 19469 2369
rect 19411 2329 19423 2363
rect 19457 2360 19469 2363
rect 50044 2360 50050 2372
rect 19457 2332 50050 2360
rect 19457 2329 19469 2332
rect 19411 2323 19469 2329
rect 50044 2320 50050 2332
rect 50102 2320 50108 2372
rect 14532 2252 14538 2304
rect 14590 2292 14596 2304
rect 50139 2295 50197 2301
rect 50139 2292 50151 2295
rect 14590 2264 50151 2292
rect 14590 2252 14596 2264
rect 50139 2261 50151 2264
rect 50185 2261 50197 2295
rect 50139 2255 50197 2261
rect 1086 2202 58862 2224
rect 1086 2150 4228 2202
rect 4280 2150 4292 2202
rect 4344 2150 4356 2202
rect 4408 2150 4420 2202
rect 4472 2150 34948 2202
rect 35000 2150 35012 2202
rect 35064 2150 35076 2202
rect 35128 2150 35140 2202
rect 35192 2150 58862 2202
rect 1086 2128 58862 2150
rect 30632 2048 30638 2100
rect 30690 2088 30696 2100
rect 31276 2088 31282 2100
rect 30690 2060 31282 2088
rect 30690 2048 30696 2060
rect 31276 2048 31282 2060
rect 31334 2048 31340 2100
rect 30172 1980 30178 2032
rect 30230 2020 30236 2032
rect 36520 2020 36526 2032
rect 30230 1992 36526 2020
rect 30230 1980 30236 1992
rect 36520 1980 36526 1992
rect 36578 1980 36584 2032
rect 29068 1844 29074 1896
rect 29126 1884 29132 1896
rect 35784 1884 35790 1896
rect 29126 1856 35790 1884
rect 29126 1844 29132 1856
rect 35784 1844 35790 1856
rect 35842 1844 35848 1896
rect 39832 1708 39838 1760
rect 39890 1748 39896 1760
rect 41304 1748 41310 1760
rect 39890 1720 41310 1748
rect 39890 1708 39896 1720
rect 41304 1708 41310 1720
rect 41362 1708 41368 1760
rect 38820 1572 38826 1624
rect 38878 1612 38884 1624
rect 39832 1612 39838 1624
rect 38878 1584 39838 1612
rect 38878 1572 38884 1584
rect 39832 1572 39838 1584
rect 39890 1572 39896 1624
rect 17936 1368 17942 1420
rect 17994 1408 18000 1420
rect 18212 1408 18218 1420
rect 17994 1380 18218 1408
rect 17994 1368 18000 1380
rect 18212 1368 18218 1380
rect 18270 1368 18276 1420
rect 19684 1368 19690 1420
rect 19742 1408 19748 1420
rect 20512 1408 20518 1420
rect 19742 1380 20518 1408
rect 19742 1368 19748 1380
rect 20512 1368 20518 1380
rect 20570 1368 20576 1420
rect 29344 1368 29350 1420
rect 29402 1408 29408 1420
rect 30264 1408 30270 1420
rect 29402 1380 30270 1408
rect 29402 1368 29408 1380
rect 30264 1368 30270 1380
rect 30322 1368 30328 1420
rect 49952 1368 49958 1420
rect 50010 1408 50016 1420
rect 50872 1408 50878 1420
rect 50010 1380 50878 1408
rect 50010 1368 50016 1380
rect 50872 1368 50878 1380
rect 50930 1368 50936 1420
rect 29160 892 29166 944
rect 29218 932 29224 944
rect 29252 932 29258 944
rect 29218 904 29258 932
rect 29218 892 29224 904
rect 29252 892 29258 904
rect 29310 892 29316 944
<< via1 >>
rect 4326 59100 4378 59152
rect 6166 59100 6218 59152
rect 45726 59100 45778 59152
rect 45910 59100 45962 59152
rect 56766 57876 56818 57928
rect 56858 57876 56910 57928
rect 34686 57808 34738 57860
rect 34870 57808 34922 57860
rect 4228 57638 4280 57690
rect 4292 57638 4344 57690
rect 4356 57638 4408 57690
rect 4420 57638 4472 57690
rect 34948 57638 35000 57690
rect 35012 57638 35064 57690
rect 35076 57638 35128 57690
rect 35140 57638 35192 57690
rect 19588 57094 19640 57146
rect 19652 57094 19704 57146
rect 19716 57094 19768 57146
rect 19780 57094 19832 57146
rect 50308 57094 50360 57146
rect 50372 57094 50424 57146
rect 50436 57094 50488 57146
rect 50500 57094 50552 57146
rect 23738 56788 23790 56840
rect 29442 56831 29494 56840
rect 29442 56797 29451 56831
rect 29451 56797 29485 56831
rect 29485 56797 29494 56831
rect 29442 56788 29494 56797
rect 39470 56720 39522 56772
rect 44898 56720 44950 56772
rect 15826 56652 15878 56704
rect 26038 56652 26090 56704
rect 4228 56550 4280 56602
rect 4292 56550 4344 56602
rect 4356 56550 4408 56602
rect 4420 56550 4472 56602
rect 34948 56550 35000 56602
rect 35012 56550 35064 56602
rect 35076 56550 35128 56602
rect 35140 56550 35192 56602
rect 646 56448 698 56500
rect 1198 56448 1250 56500
rect 1750 56448 1802 56500
rect 2670 56448 2722 56500
rect 13618 56448 13670 56500
rect 186 56380 238 56432
rect 1290 56380 1342 56432
rect 14446 56380 14498 56432
rect 21070 56380 21122 56432
rect 23738 56448 23790 56500
rect 28062 56380 28114 56432
rect 28154 56380 28206 56432
rect 31190 56380 31242 56432
rect 31926 56448 31978 56500
rect 35974 56448 36026 56500
rect 36066 56448 36118 56500
rect 41402 56448 41454 56500
rect 41494 56448 41546 56500
rect 54834 56448 54886 56500
rect 40114 56380 40166 56432
rect 40206 56380 40258 56432
rect 10858 56312 10910 56364
rect 26682 56312 26734 56364
rect 26774 56312 26826 56364
rect 35882 56312 35934 56364
rect 35974 56312 36026 56364
rect 10582 56244 10634 56296
rect 15918 56244 15970 56296
rect 19966 56244 20018 56296
rect 24014 56244 24066 56296
rect 29442 56244 29494 56296
rect 29718 56244 29770 56296
rect 32938 56244 32990 56296
rect 33030 56244 33082 56296
rect 36066 56244 36118 56296
rect 36526 56312 36578 56364
rect 41126 56312 41178 56364
rect 41310 56380 41362 56432
rect 51154 56380 51206 56432
rect 52718 56312 52770 56364
rect 40666 56244 40718 56296
rect 40758 56244 40810 56296
rect 57502 56244 57554 56296
rect 4050 56176 4102 56228
rect 16470 56176 16522 56228
rect 21622 56176 21674 56228
rect 26866 56176 26918 56228
rect 27050 56176 27102 56228
rect 31558 56176 31610 56228
rect 31650 56176 31702 56228
rect 33030 56108 33082 56160
rect 33214 56176 33266 56228
rect 41402 56108 41454 56160
rect 41586 56176 41638 56228
rect 43242 56176 43294 56228
rect 44162 56176 44214 56228
rect 45358 56176 45410 56228
rect 45450 56176 45502 56228
rect 48578 56176 48630 56228
rect 41678 56108 41730 56160
rect 44898 56108 44950 56160
rect 55938 56108 55990 56160
rect 19588 56006 19640 56058
rect 19652 56006 19704 56058
rect 19716 56006 19768 56058
rect 19780 56006 19832 56058
rect 50308 56006 50360 56058
rect 50372 56006 50424 56058
rect 50436 56006 50488 56058
rect 50500 56006 50552 56058
rect 9846 55904 9898 55956
rect 29810 55904 29862 55956
rect 31650 55904 31702 55956
rect 31742 55904 31794 55956
rect 33214 55904 33266 55956
rect 35422 55904 35474 55956
rect 38642 55904 38694 55956
rect 39654 55904 39706 55956
rect 58054 55904 58106 55956
rect 8098 55836 8150 55888
rect 44162 55836 44214 55888
rect 44714 55836 44766 55888
rect 59066 55836 59118 55888
rect 8558 55768 8610 55820
rect 13066 55768 13118 55820
rect 20150 55768 20202 55820
rect 26222 55768 26274 55820
rect 37538 55768 37590 55820
rect 37630 55768 37682 55820
rect 40574 55768 40626 55820
rect 40666 55768 40718 55820
rect 59618 55768 59670 55820
rect 7270 55700 7322 55752
rect 18034 55700 18086 55752
rect 19414 55700 19466 55752
rect 26774 55700 26826 55752
rect 26866 55700 26918 55752
rect 33858 55700 33910 55752
rect 33950 55700 34002 55752
rect 10490 55632 10542 55684
rect 17482 55632 17534 55684
rect 18678 55632 18730 55684
rect 22726 55632 22778 55684
rect 26222 55632 26274 55684
rect 27510 55632 27562 55684
rect 31926 55632 31978 55684
rect 32018 55632 32070 55684
rect 35330 55632 35382 55684
rect 35882 55700 35934 55752
rect 38550 55700 38602 55752
rect 38642 55700 38694 55752
rect 53270 55700 53322 55752
rect 37078 55632 37130 55684
rect 38090 55632 38142 55684
rect 42230 55632 42282 55684
rect 44622 55632 44674 55684
rect 54374 55632 54426 55684
rect 13250 55564 13302 55616
rect 20978 55564 21030 55616
rect 21070 55564 21122 55616
rect 23278 55564 23330 55616
rect 25946 55564 25998 55616
rect 27418 55564 27470 55616
rect 27602 55564 27654 55616
rect 31098 55564 31150 55616
rect 31190 55564 31242 55616
rect 38274 55564 38326 55616
rect 41402 55564 41454 55616
rect 41494 55564 41546 55616
rect 47014 55564 47066 55616
rect 52442 55607 52494 55616
rect 52442 55573 52451 55607
rect 52451 55573 52485 55607
rect 52485 55573 52494 55607
rect 52442 55564 52494 55573
rect 4228 55462 4280 55514
rect 4292 55462 4344 55514
rect 4356 55462 4408 55514
rect 4420 55462 4472 55514
rect 34948 55462 35000 55514
rect 35012 55462 35064 55514
rect 35076 55462 35128 55514
rect 35140 55462 35192 55514
rect 17574 55360 17626 55412
rect 20702 55360 20754 55412
rect 23370 55360 23422 55412
rect 30914 55360 30966 55412
rect 4878 55292 4930 55344
rect 6258 55292 6310 55344
rect 6442 55292 6494 55344
rect 8190 55292 8242 55344
rect 14998 55292 15050 55344
rect 17022 55292 17074 55344
rect 20058 55292 20110 55344
rect 2762 55224 2814 55276
rect 3958 55224 4010 55276
rect 5890 55224 5942 55276
rect 6810 55224 6862 55276
rect 6994 55224 7046 55276
rect 8006 55224 8058 55276
rect 8282 55224 8334 55276
rect 9570 55224 9622 55276
rect 11686 55224 11738 55276
rect 12146 55224 12198 55276
rect 13802 55224 13854 55276
rect 15090 55224 15142 55276
rect 18586 55224 18638 55276
rect 19138 55224 19190 55276
rect 19874 55224 19926 55276
rect 20610 55224 20662 55276
rect 20978 55292 21030 55344
rect 24014 55292 24066 55344
rect 29074 55292 29126 55344
rect 30270 55292 30322 55344
rect 24842 55224 24894 55276
rect 26038 55224 26090 55276
rect 28246 55224 28298 55276
rect 29626 55224 29678 55276
rect 31466 55360 31518 55412
rect 31834 55360 31886 55412
rect 31098 55292 31150 55344
rect 32018 55292 32070 55344
rect 32754 55292 32806 55344
rect 32938 55360 32990 55412
rect 36986 55360 37038 55412
rect 37078 55360 37130 55412
rect 41310 55360 41362 55412
rect 41678 55360 41730 55412
rect 43794 55360 43846 55412
rect 43886 55360 43938 55412
rect 46462 55360 46514 55412
rect 39470 55292 39522 55344
rect 43610 55292 43662 55344
rect 50142 55292 50194 55344
rect 31006 55156 31058 55208
rect 32202 55224 32254 55276
rect 33030 55224 33082 55276
rect 32386 55156 32438 55208
rect 33950 55224 34002 55276
rect 33214 55156 33266 55208
rect 30914 55088 30966 55140
rect 32938 55088 32990 55140
rect 35330 55224 35382 55276
rect 41310 55224 41362 55276
rect 41494 55224 41546 55276
rect 51706 55224 51758 55276
rect 43886 55088 43938 55140
rect 33858 55020 33910 55072
rect 37630 55020 37682 55072
rect 19588 54918 19640 54970
rect 19652 54918 19704 54970
rect 19716 54918 19768 54970
rect 19780 54918 19832 54970
rect 50308 54918 50360 54970
rect 50372 54918 50424 54970
rect 50436 54918 50488 54970
rect 50500 54918 50552 54970
rect 4050 54476 4102 54528
rect 19322 54544 19374 54596
rect 18126 54519 18178 54528
rect 18126 54485 18135 54519
rect 18135 54485 18169 54519
rect 18169 54485 18178 54519
rect 18126 54476 18178 54485
rect 22542 54476 22594 54528
rect 23554 54476 23606 54528
rect 4228 54374 4280 54426
rect 4292 54374 4344 54426
rect 4356 54374 4408 54426
rect 4420 54374 4472 54426
rect 34948 54374 35000 54426
rect 35012 54374 35064 54426
rect 35076 54374 35128 54426
rect 35140 54374 35192 54426
rect 22542 54272 22594 54324
rect 48946 54272 48998 54324
rect 21714 54204 21766 54256
rect 27142 54204 27194 54256
rect 22726 54068 22778 54120
rect 19588 53830 19640 53882
rect 19652 53830 19704 53882
rect 19716 53830 19768 53882
rect 19780 53830 19832 53882
rect 50308 53830 50360 53882
rect 50372 53830 50424 53882
rect 50436 53830 50488 53882
rect 50500 53830 50552 53882
rect 30638 53728 30690 53780
rect 4228 53286 4280 53338
rect 4292 53286 4344 53338
rect 4356 53286 4408 53338
rect 4420 53286 4472 53338
rect 34948 53286 35000 53338
rect 35012 53286 35064 53338
rect 35076 53286 35128 53338
rect 35140 53286 35192 53338
rect 23370 53184 23422 53236
rect 39010 53048 39062 53100
rect 39562 53048 39614 53100
rect 12330 52980 12382 53032
rect 19588 52742 19640 52794
rect 19652 52742 19704 52794
rect 19716 52742 19768 52794
rect 19780 52742 19832 52794
rect 50308 52742 50360 52794
rect 50372 52742 50424 52794
rect 50436 52742 50488 52794
rect 50500 52742 50552 52794
rect 5062 52368 5114 52420
rect 35882 52368 35934 52420
rect 7638 52343 7690 52352
rect 7638 52309 7647 52343
rect 7647 52309 7681 52343
rect 7681 52309 7690 52343
rect 7638 52300 7690 52309
rect 39654 52343 39706 52352
rect 39654 52309 39663 52343
rect 39663 52309 39697 52343
rect 39697 52309 39706 52343
rect 39654 52300 39706 52309
rect 4228 52198 4280 52250
rect 4292 52198 4344 52250
rect 4356 52198 4408 52250
rect 4420 52198 4472 52250
rect 34948 52198 35000 52250
rect 35012 52198 35064 52250
rect 35076 52198 35128 52250
rect 35140 52198 35192 52250
rect 19588 51654 19640 51706
rect 19652 51654 19704 51706
rect 19716 51654 19768 51706
rect 19780 51654 19832 51706
rect 50308 51654 50360 51706
rect 50372 51654 50424 51706
rect 50436 51654 50488 51706
rect 50500 51654 50552 51706
rect 10858 51459 10910 51468
rect 10858 51425 10867 51459
rect 10867 51425 10901 51459
rect 10901 51425 10910 51459
rect 10858 51416 10910 51425
rect 4228 51110 4280 51162
rect 4292 51110 4344 51162
rect 4356 51110 4408 51162
rect 4420 51110 4472 51162
rect 34948 51110 35000 51162
rect 35012 51110 35064 51162
rect 35076 51110 35128 51162
rect 35140 51110 35192 51162
rect 13802 51008 13854 51060
rect 14906 51008 14958 51060
rect 18218 50847 18270 50856
rect 18218 50813 18227 50847
rect 18227 50813 18261 50847
rect 18261 50813 18270 50847
rect 18218 50804 18270 50813
rect 28890 50847 28942 50856
rect 28890 50813 28899 50847
rect 28899 50813 28933 50847
rect 28933 50813 28942 50847
rect 28890 50804 28942 50813
rect 19588 50566 19640 50618
rect 19652 50566 19704 50618
rect 19716 50566 19768 50618
rect 19780 50566 19832 50618
rect 50308 50566 50360 50618
rect 50372 50566 50424 50618
rect 50436 50566 50488 50618
rect 50500 50566 50552 50618
rect 4228 50022 4280 50074
rect 4292 50022 4344 50074
rect 4356 50022 4408 50074
rect 4420 50022 4472 50074
rect 34948 50022 35000 50074
rect 35012 50022 35064 50074
rect 35076 50022 35128 50074
rect 35140 50022 35192 50074
rect 16470 49716 16522 49768
rect 19588 49478 19640 49530
rect 19652 49478 19704 49530
rect 19716 49478 19768 49530
rect 19780 49478 19832 49530
rect 50308 49478 50360 49530
rect 50372 49478 50424 49530
rect 50436 49478 50488 49530
rect 50500 49478 50552 49530
rect 18862 49036 18914 49088
rect 4228 48934 4280 48986
rect 4292 48934 4344 48986
rect 4356 48934 4408 48986
rect 4420 48934 4472 48986
rect 34948 48934 35000 48986
rect 35012 48934 35064 48986
rect 35076 48934 35128 48986
rect 35140 48934 35192 48986
rect 13710 48628 13762 48680
rect 34042 48671 34094 48680
rect 34042 48637 34051 48671
rect 34051 48637 34085 48671
rect 34085 48637 34094 48671
rect 34042 48628 34094 48637
rect 19588 48390 19640 48442
rect 19652 48390 19704 48442
rect 19716 48390 19768 48442
rect 19780 48390 19832 48442
rect 50308 48390 50360 48442
rect 50372 48390 50424 48442
rect 50436 48390 50488 48442
rect 50500 48390 50552 48442
rect 8650 48288 8702 48340
rect 8742 48288 8794 48340
rect 18862 48288 18914 48340
rect 18954 48288 19006 48340
rect 24198 48288 24250 48340
rect 26406 48288 26458 48340
rect 29350 48288 29402 48340
rect 30178 48288 30230 48340
rect 34594 48288 34646 48340
rect 34686 48288 34738 48340
rect 37998 48288 38050 48340
rect 38090 48288 38142 48340
rect 35422 48220 35474 48272
rect 51154 48220 51206 48272
rect 51246 48220 51298 48272
rect 35514 48152 35566 48204
rect 34410 47948 34462 48000
rect 4228 47846 4280 47898
rect 4292 47846 4344 47898
rect 4356 47846 4408 47898
rect 4420 47846 4472 47898
rect 34948 47846 35000 47898
rect 35012 47846 35064 47898
rect 35076 47846 35128 47898
rect 35140 47846 35192 47898
rect 19588 47302 19640 47354
rect 19652 47302 19704 47354
rect 19716 47302 19768 47354
rect 19780 47302 19832 47354
rect 50308 47302 50360 47354
rect 50372 47302 50424 47354
rect 50436 47302 50488 47354
rect 50500 47302 50552 47354
rect 26866 46996 26918 47048
rect 10306 46928 10358 46980
rect 10582 46928 10634 46980
rect 17206 46928 17258 46980
rect 17574 46928 17626 46980
rect 26590 46928 26642 46980
rect 27142 46928 27194 46980
rect 4228 46758 4280 46810
rect 4292 46758 4344 46810
rect 4356 46758 4408 46810
rect 4420 46758 4472 46810
rect 34948 46758 35000 46810
rect 35012 46758 35064 46810
rect 35076 46758 35128 46810
rect 35140 46758 35192 46810
rect 20518 46452 20570 46504
rect 55110 46452 55162 46504
rect 5430 46316 5482 46368
rect 19588 46214 19640 46266
rect 19652 46214 19704 46266
rect 19716 46214 19768 46266
rect 19780 46214 19832 46266
rect 50308 46214 50360 46266
rect 50372 46214 50424 46266
rect 50436 46214 50488 46266
rect 50500 46214 50552 46266
rect 25946 46112 25998 46164
rect 26130 46112 26182 46164
rect 21346 45840 21398 45892
rect 9202 45815 9254 45824
rect 9202 45781 9211 45815
rect 9211 45781 9245 45815
rect 9245 45781 9254 45815
rect 9202 45772 9254 45781
rect 20518 45815 20570 45824
rect 20518 45781 20527 45815
rect 20527 45781 20561 45815
rect 20561 45781 20570 45815
rect 20518 45772 20570 45781
rect 23186 45772 23238 45824
rect 4228 45670 4280 45722
rect 4292 45670 4344 45722
rect 4356 45670 4408 45722
rect 4420 45670 4472 45722
rect 34948 45670 35000 45722
rect 35012 45670 35064 45722
rect 35076 45670 35128 45722
rect 35140 45670 35192 45722
rect 7454 45568 7506 45620
rect 7730 45568 7782 45620
rect 7914 45568 7966 45620
rect 20518 45568 20570 45620
rect 26222 45500 26274 45552
rect 26590 45500 26642 45552
rect 38826 45500 38878 45552
rect 39010 45500 39062 45552
rect 9570 45364 9622 45416
rect 29442 45407 29494 45416
rect 29442 45373 29451 45407
rect 29451 45373 29485 45407
rect 29485 45373 29494 45407
rect 29442 45364 29494 45373
rect 17850 45296 17902 45348
rect 19588 45126 19640 45178
rect 19652 45126 19704 45178
rect 19716 45126 19768 45178
rect 19780 45126 19832 45178
rect 50308 45126 50360 45178
rect 50372 45126 50424 45178
rect 50436 45126 50488 45178
rect 50500 45126 50552 45178
rect 16378 44684 16430 44736
rect 4228 44582 4280 44634
rect 4292 44582 4344 44634
rect 4356 44582 4408 44634
rect 4420 44582 4472 44634
rect 34948 44582 35000 44634
rect 35012 44582 35064 44634
rect 35076 44582 35128 44634
rect 35140 44582 35192 44634
rect 26866 44344 26918 44396
rect 5154 44208 5206 44260
rect 29902 44276 29954 44328
rect 36618 44319 36670 44328
rect 36618 44285 36627 44319
rect 36627 44285 36661 44319
rect 36661 44285 36670 44319
rect 36618 44276 36670 44285
rect 38182 44319 38234 44328
rect 38182 44285 38191 44319
rect 38191 44285 38225 44319
rect 38225 44285 38234 44319
rect 38182 44276 38234 44285
rect 45542 44140 45594 44192
rect 45726 44140 45778 44192
rect 19588 44038 19640 44090
rect 19652 44038 19704 44090
rect 19716 44038 19768 44090
rect 19780 44038 19832 44090
rect 50308 44038 50360 44090
rect 50372 44038 50424 44090
rect 50436 44038 50488 44090
rect 50500 44038 50552 44090
rect 44898 43979 44950 43988
rect 44898 43945 44907 43979
rect 44907 43945 44941 43979
rect 44941 43945 44950 43979
rect 44898 43936 44950 43945
rect 48302 43936 48354 43988
rect 48302 43800 48354 43852
rect 37446 43775 37498 43784
rect 37446 43741 37455 43775
rect 37455 43741 37489 43775
rect 37489 43741 37498 43775
rect 37446 43732 37498 43741
rect 30270 43664 30322 43716
rect 50970 43732 51022 43784
rect 51062 43732 51114 43784
rect 20058 43596 20110 43648
rect 23370 43596 23422 43648
rect 4228 43494 4280 43546
rect 4292 43494 4344 43546
rect 4356 43494 4408 43546
rect 4420 43494 4472 43546
rect 34948 43494 35000 43546
rect 35012 43494 35064 43546
rect 35076 43494 35128 43546
rect 35140 43494 35192 43546
rect 14998 43435 15050 43444
rect 14998 43401 15007 43435
rect 15007 43401 15041 43435
rect 15041 43401 15050 43435
rect 14998 43392 15050 43401
rect 34594 43324 34646 43376
rect 34778 43324 34830 43376
rect 20150 43120 20202 43172
rect 33858 43052 33910 43104
rect 19588 42950 19640 43002
rect 19652 42950 19704 43002
rect 19716 42950 19768 43002
rect 19780 42950 19832 43002
rect 50308 42950 50360 43002
rect 50372 42950 50424 43002
rect 50436 42950 50488 43002
rect 50500 42950 50552 43002
rect 4228 42406 4280 42458
rect 4292 42406 4344 42458
rect 4356 42406 4408 42458
rect 4420 42406 4472 42458
rect 34948 42406 35000 42458
rect 35012 42406 35064 42458
rect 35076 42406 35128 42458
rect 35140 42406 35192 42458
rect 9938 42211 9990 42220
rect 9938 42177 9947 42211
rect 9947 42177 9981 42211
rect 9981 42177 9990 42211
rect 9938 42168 9990 42177
rect 13526 42100 13578 42152
rect 19588 41862 19640 41914
rect 19652 41862 19704 41914
rect 19716 41862 19768 41914
rect 19780 41862 19832 41914
rect 50308 41862 50360 41914
rect 50372 41862 50424 41914
rect 50436 41862 50488 41914
rect 50500 41862 50552 41914
rect 4228 41318 4280 41370
rect 4292 41318 4344 41370
rect 4356 41318 4408 41370
rect 4420 41318 4472 41370
rect 34948 41318 35000 41370
rect 35012 41318 35064 41370
rect 35076 41318 35128 41370
rect 35140 41318 35192 41370
rect 19966 41259 20018 41268
rect 19966 41225 19975 41259
rect 19975 41225 20009 41259
rect 20009 41225 20018 41259
rect 19966 41216 20018 41225
rect 28338 41012 28390 41064
rect 24198 40944 24250 40996
rect 19588 40774 19640 40826
rect 19652 40774 19704 40826
rect 19716 40774 19768 40826
rect 19780 40774 19832 40826
rect 50308 40774 50360 40826
rect 50372 40774 50424 40826
rect 50436 40774 50488 40826
rect 50500 40774 50552 40826
rect 27142 40332 27194 40384
rect 50970 40332 51022 40384
rect 4228 40230 4280 40282
rect 4292 40230 4344 40282
rect 4356 40230 4408 40282
rect 4420 40230 4472 40282
rect 34948 40230 35000 40282
rect 35012 40230 35064 40282
rect 35076 40230 35128 40282
rect 35140 40230 35192 40282
rect 4970 40103 5022 40112
rect 4970 40069 4979 40103
rect 4979 40069 5013 40103
rect 5013 40069 5022 40103
rect 4970 40060 5022 40069
rect 14630 40103 14682 40112
rect 14630 40069 14639 40103
rect 14639 40069 14673 40103
rect 14673 40069 14682 40103
rect 14630 40060 14682 40069
rect 28798 40060 28850 40112
rect 19588 39686 19640 39738
rect 19652 39686 19704 39738
rect 19716 39686 19768 39738
rect 19780 39686 19832 39738
rect 50308 39686 50360 39738
rect 50372 39686 50424 39738
rect 50436 39686 50488 39738
rect 50500 39686 50552 39738
rect 20518 39380 20570 39432
rect 23370 39380 23422 39432
rect 27510 39380 27562 39432
rect 7362 39312 7414 39364
rect 7546 39312 7598 39364
rect 5246 39244 5298 39296
rect 36986 39287 37038 39296
rect 36986 39253 36995 39287
rect 36995 39253 37029 39287
rect 37029 39253 37038 39287
rect 36986 39244 37038 39253
rect 49590 39244 49642 39296
rect 4228 39142 4280 39194
rect 4292 39142 4344 39194
rect 4356 39142 4408 39194
rect 4420 39142 4472 39194
rect 34948 39142 35000 39194
rect 35012 39142 35064 39194
rect 35076 39142 35128 39194
rect 35140 39142 35192 39194
rect 19138 39040 19190 39092
rect 19588 38598 19640 38650
rect 19652 38598 19704 38650
rect 19716 38598 19768 38650
rect 19780 38598 19832 38650
rect 50308 38598 50360 38650
rect 50372 38598 50424 38650
rect 50436 38598 50488 38650
rect 50500 38598 50552 38650
rect 28982 38156 29034 38208
rect 4228 38054 4280 38106
rect 4292 38054 4344 38106
rect 4356 38054 4408 38106
rect 4420 38054 4472 38106
rect 34948 38054 35000 38106
rect 35012 38054 35064 38106
rect 35076 38054 35128 38106
rect 35140 38054 35192 38106
rect 19588 37510 19640 37562
rect 19652 37510 19704 37562
rect 19716 37510 19768 37562
rect 19780 37510 19832 37562
rect 50308 37510 50360 37562
rect 50372 37510 50424 37562
rect 50436 37510 50488 37562
rect 50500 37510 50552 37562
rect 21806 37451 21858 37460
rect 21806 37417 21815 37451
rect 21815 37417 21849 37451
rect 21849 37417 21858 37451
rect 21806 37408 21858 37417
rect 8650 37272 8702 37324
rect 8742 37272 8794 37324
rect 29902 37272 29954 37324
rect 29994 37272 30046 37324
rect 37446 37272 37498 37324
rect 46278 37272 46330 37324
rect 6810 37204 6862 37256
rect 1106 37068 1158 37120
rect 11134 37111 11186 37120
rect 11134 37077 11143 37111
rect 11143 37077 11177 37111
rect 11177 37077 11186 37111
rect 11134 37068 11186 37077
rect 38550 37068 38602 37120
rect 4228 36966 4280 37018
rect 4292 36966 4344 37018
rect 4356 36966 4408 37018
rect 4420 36966 4472 37018
rect 34948 36966 35000 37018
rect 35012 36966 35064 37018
rect 35076 36966 35128 37018
rect 35140 36966 35192 37018
rect 19414 36907 19466 36916
rect 19414 36873 19423 36907
rect 19423 36873 19457 36907
rect 19457 36873 19466 36907
rect 19414 36864 19466 36873
rect 34318 36728 34370 36780
rect 3774 36660 3826 36712
rect 11778 36703 11830 36712
rect 11778 36669 11787 36703
rect 11787 36669 11821 36703
rect 11821 36669 11830 36703
rect 11778 36660 11830 36669
rect 35238 36660 35290 36712
rect 40758 36592 40810 36644
rect 19588 36422 19640 36474
rect 19652 36422 19704 36474
rect 19716 36422 19768 36474
rect 19780 36422 19832 36474
rect 50308 36422 50360 36474
rect 50372 36422 50424 36474
rect 50436 36422 50488 36474
rect 50500 36422 50552 36474
rect 25946 36320 25998 36372
rect 26130 36320 26182 36372
rect 6350 36023 6402 36032
rect 6350 35989 6359 36023
rect 6359 35989 6393 36023
rect 6393 35989 6402 36023
rect 6350 35980 6402 35989
rect 26222 35980 26274 36032
rect 26406 35980 26458 36032
rect 38090 36023 38142 36032
rect 38090 35989 38099 36023
rect 38099 35989 38133 36023
rect 38133 35989 38142 36023
rect 38090 35980 38142 35989
rect 4228 35878 4280 35930
rect 4292 35878 4344 35930
rect 4356 35878 4408 35930
rect 4420 35878 4472 35930
rect 34948 35878 35000 35930
rect 35012 35878 35064 35930
rect 35076 35878 35128 35930
rect 35140 35878 35192 35930
rect 38366 35819 38418 35828
rect 38366 35785 38375 35819
rect 38375 35785 38409 35819
rect 38409 35785 38418 35819
rect 38366 35776 38418 35785
rect 21438 35572 21490 35624
rect 55662 35615 55714 35624
rect 55662 35581 55671 35615
rect 55671 35581 55705 35615
rect 55705 35581 55714 35615
rect 55662 35572 55714 35581
rect 19588 35334 19640 35386
rect 19652 35334 19704 35386
rect 19716 35334 19768 35386
rect 19780 35334 19832 35386
rect 50308 35334 50360 35386
rect 50372 35334 50424 35386
rect 50436 35334 50488 35386
rect 50500 35334 50552 35386
rect 1106 34892 1158 34944
rect 4228 34790 4280 34842
rect 4292 34790 4344 34842
rect 4356 34790 4408 34842
rect 4420 34790 4472 34842
rect 34948 34790 35000 34842
rect 35012 34790 35064 34842
rect 35076 34790 35128 34842
rect 35140 34790 35192 34842
rect 7362 34484 7414 34536
rect 7638 34484 7690 34536
rect 23002 34484 23054 34536
rect 23186 34484 23238 34536
rect 44990 34484 45042 34536
rect 19588 34246 19640 34298
rect 19652 34246 19704 34298
rect 19716 34246 19768 34298
rect 19780 34246 19832 34298
rect 50308 34246 50360 34298
rect 50372 34246 50424 34298
rect 50436 34246 50488 34298
rect 50500 34246 50552 34298
rect 42046 33804 42098 33856
rect 48486 33804 48538 33856
rect 48670 33804 48722 33856
rect 4228 33702 4280 33754
rect 4292 33702 4344 33754
rect 4356 33702 4408 33754
rect 4420 33702 4472 33754
rect 34948 33702 35000 33754
rect 35012 33702 35064 33754
rect 35076 33702 35128 33754
rect 35140 33702 35192 33754
rect 19588 33158 19640 33210
rect 19652 33158 19704 33210
rect 19716 33158 19768 33210
rect 19780 33158 19832 33210
rect 50308 33158 50360 33210
rect 50372 33158 50424 33210
rect 50436 33158 50488 33210
rect 50500 33158 50552 33210
rect 22634 32920 22686 32972
rect 9202 32716 9254 32768
rect 9478 32716 9530 32768
rect 11870 32759 11922 32768
rect 11870 32725 11879 32759
rect 11879 32725 11913 32759
rect 11913 32725 11922 32759
rect 11870 32716 11922 32725
rect 22634 32716 22686 32768
rect 32478 32716 32530 32768
rect 4228 32614 4280 32666
rect 4292 32614 4344 32666
rect 4356 32614 4408 32666
rect 4420 32614 4472 32666
rect 34948 32614 35000 32666
rect 35012 32614 35064 32666
rect 35076 32614 35128 32666
rect 35140 32614 35192 32666
rect 2486 32512 2538 32564
rect 11870 32512 11922 32564
rect 23186 32444 23238 32496
rect 23554 32444 23606 32496
rect 8742 32376 8794 32428
rect 9202 32376 9254 32428
rect 26958 32376 27010 32428
rect 27142 32376 27194 32428
rect 19588 32070 19640 32122
rect 19652 32070 19704 32122
rect 19716 32070 19768 32122
rect 19780 32070 19832 32122
rect 50308 32070 50360 32122
rect 50372 32070 50424 32122
rect 50436 32070 50488 32122
rect 50500 32070 50552 32122
rect 21990 31764 22042 31816
rect 4228 31526 4280 31578
rect 4292 31526 4344 31578
rect 4356 31526 4408 31578
rect 4420 31526 4472 31578
rect 34948 31526 35000 31578
rect 35012 31526 35064 31578
rect 35076 31526 35128 31578
rect 35140 31526 35192 31578
rect 8742 31220 8794 31272
rect 11042 31220 11094 31272
rect 11226 31263 11278 31272
rect 11226 31229 11235 31263
rect 11235 31229 11269 31263
rect 11269 31229 11278 31263
rect 11226 31220 11278 31229
rect 38826 31220 38878 31272
rect 8834 31084 8886 31136
rect 9018 31084 9070 31136
rect 28430 31084 28482 31136
rect 19588 30982 19640 31034
rect 19652 30982 19704 31034
rect 19716 30982 19768 31034
rect 19780 30982 19832 31034
rect 50308 30982 50360 31034
rect 50372 30982 50424 31034
rect 50436 30982 50488 31034
rect 50500 30982 50552 31034
rect 11042 30880 11094 30932
rect 27878 30880 27930 30932
rect 8742 30812 8794 30864
rect 28706 30812 28758 30864
rect 4228 30438 4280 30490
rect 4292 30438 4344 30490
rect 4356 30438 4408 30490
rect 4420 30438 4472 30490
rect 34948 30438 35000 30490
rect 35012 30438 35064 30490
rect 35076 30438 35128 30490
rect 35140 30438 35192 30490
rect 8466 30132 8518 30184
rect 13158 30132 13210 30184
rect 14998 30132 15050 30184
rect 29534 30132 29586 30184
rect 48118 30175 48170 30184
rect 48118 30141 48127 30175
rect 48127 30141 48161 30175
rect 48161 30141 48170 30175
rect 48118 30132 48170 30141
rect 48486 30175 48538 30184
rect 48486 30141 48495 30175
rect 48495 30141 48529 30175
rect 48529 30141 48538 30175
rect 48486 30132 48538 30141
rect 39930 30064 39982 30116
rect 8834 29996 8886 30048
rect 9018 29996 9070 30048
rect 25486 29996 25538 30048
rect 19588 29894 19640 29946
rect 19652 29894 19704 29946
rect 19716 29894 19768 29946
rect 19780 29894 19832 29946
rect 50308 29894 50360 29946
rect 50372 29894 50424 29946
rect 50436 29894 50488 29946
rect 50500 29894 50552 29946
rect 13158 29792 13210 29844
rect 27234 29792 27286 29844
rect 1014 29724 1066 29776
rect 48486 29724 48538 29776
rect 7730 29656 7782 29708
rect 48118 29656 48170 29708
rect 8466 29588 8518 29640
rect 27694 29588 27746 29640
rect 8834 29520 8886 29572
rect 25854 29520 25906 29572
rect 15642 29495 15694 29504
rect 15642 29461 15651 29495
rect 15651 29461 15685 29495
rect 15685 29461 15694 29495
rect 15642 29452 15694 29461
rect 4228 29350 4280 29402
rect 4292 29350 4344 29402
rect 4356 29350 4408 29402
rect 4420 29350 4472 29402
rect 34948 29350 35000 29402
rect 35012 29350 35064 29402
rect 35076 29350 35128 29402
rect 35140 29350 35192 29402
rect 27142 29248 27194 29300
rect 8834 29112 8886 29164
rect 26314 29112 26366 29164
rect 12054 29044 12106 29096
rect 19046 28976 19098 29028
rect 19138 28976 19190 29028
rect 24014 28976 24066 29028
rect 24106 28976 24158 29028
rect 34686 28976 34738 29028
rect 34778 28976 34830 29028
rect 48302 28976 48354 29028
rect 48670 28976 48722 29028
rect 24382 28908 24434 28960
rect 19588 28806 19640 28858
rect 19652 28806 19704 28858
rect 19716 28806 19768 28858
rect 19780 28806 19832 28858
rect 50308 28806 50360 28858
rect 50372 28806 50424 28858
rect 50436 28806 50488 28858
rect 50500 28806 50552 28858
rect 27602 28747 27654 28756
rect 27602 28713 27611 28747
rect 27611 28713 27645 28747
rect 27645 28713 27654 28747
rect 27602 28704 27654 28713
rect 23278 28636 23330 28688
rect 23462 28636 23514 28688
rect 3682 28364 3734 28416
rect 34778 28407 34830 28416
rect 34778 28373 34787 28407
rect 34787 28373 34821 28407
rect 34821 28373 34830 28407
rect 34778 28364 34830 28373
rect 4228 28262 4280 28314
rect 4292 28262 4344 28314
rect 4356 28262 4408 28314
rect 4420 28262 4472 28314
rect 34948 28262 35000 28314
rect 35012 28262 35064 28314
rect 35076 28262 35128 28314
rect 35140 28262 35192 28314
rect 13894 28160 13946 28212
rect 34778 28160 34830 28212
rect 8558 28024 8610 28076
rect 8926 28024 8978 28076
rect 25394 28024 25446 28076
rect 8834 27956 8886 28008
rect 24290 27956 24342 28008
rect 37814 27999 37866 28008
rect 37814 27965 37823 27999
rect 37823 27965 37857 27999
rect 37857 27965 37866 27999
rect 37814 27956 37866 27965
rect 8558 27820 8610 27872
rect 22818 27820 22870 27872
rect 19588 27718 19640 27770
rect 19652 27718 19704 27770
rect 19716 27718 19768 27770
rect 19780 27718 19832 27770
rect 50308 27718 50360 27770
rect 50372 27718 50424 27770
rect 50436 27718 50488 27770
rect 50500 27718 50552 27770
rect 9294 27616 9346 27668
rect 9478 27616 9530 27668
rect 13342 27616 13394 27668
rect 13894 27616 13946 27668
rect 26406 27616 26458 27668
rect 26498 27616 26550 27668
rect 28430 27616 28482 27668
rect 29166 27616 29218 27668
rect 18862 27548 18914 27600
rect 18954 27548 19006 27600
rect 4228 27174 4280 27226
rect 4292 27174 4344 27226
rect 4356 27174 4408 27226
rect 4420 27174 4472 27226
rect 34948 27174 35000 27226
rect 35012 27174 35064 27226
rect 35076 27174 35128 27226
rect 35140 27174 35192 27226
rect 8420 26970 8472 27022
rect 8834 27004 8886 27056
rect 16562 27004 16614 27056
rect 8558 26868 8610 26920
rect 8834 26868 8886 26920
rect 20702 26868 20754 26920
rect 25946 26868 25998 26920
rect 26130 26868 26182 26920
rect 16562 26800 16614 26852
rect 23002 26800 23054 26852
rect 24658 26800 24710 26852
rect 7822 26732 7874 26784
rect 8190 26732 8242 26784
rect 8696 26732 8748 26784
rect 29626 26732 29678 26784
rect 19588 26630 19640 26682
rect 19652 26630 19704 26682
rect 19716 26630 19768 26682
rect 19780 26630 19832 26682
rect 50308 26630 50360 26682
rect 50372 26630 50424 26682
rect 50436 26630 50488 26682
rect 50500 26630 50552 26682
rect 8696 26528 8748 26580
rect 22910 26528 22962 26580
rect 6810 26392 6862 26444
rect 12146 26324 12198 26376
rect 32938 26324 32990 26376
rect 25026 26299 25078 26308
rect 25026 26265 25035 26299
rect 25035 26265 25069 26299
rect 25069 26265 25078 26299
rect 25026 26256 25078 26265
rect 31650 26256 31702 26308
rect 38734 26188 38786 26240
rect 39010 26188 39062 26240
rect 4228 26086 4280 26138
rect 4292 26086 4344 26138
rect 4356 26086 4408 26138
rect 4420 26086 4472 26138
rect 34948 26086 35000 26138
rect 35012 26086 35064 26138
rect 35076 26086 35128 26138
rect 35140 26086 35192 26138
rect 13618 26027 13670 26036
rect 13618 25993 13627 26027
rect 13627 25993 13661 26027
rect 13661 25993 13670 26027
rect 13618 25984 13670 25993
rect 8558 25780 8610 25832
rect 20334 25848 20386 25900
rect 37630 25780 37682 25832
rect 20334 25712 20386 25764
rect 20426 25712 20478 25764
rect 8190 25644 8242 25696
rect 8696 25644 8748 25696
rect 8834 25644 8886 25696
rect 22450 25644 22502 25696
rect 19588 25542 19640 25594
rect 19652 25542 19704 25594
rect 19716 25542 19768 25594
rect 19780 25542 19832 25594
rect 50308 25542 50360 25594
rect 50372 25542 50424 25594
rect 50436 25542 50488 25594
rect 50500 25542 50552 25594
rect 8190 25440 8242 25492
rect 22634 25440 22686 25492
rect 8696 25372 8748 25424
rect 21622 25372 21674 25424
rect 37630 25236 37682 25288
rect 44806 25236 44858 25288
rect 31558 25100 31610 25152
rect 4228 24998 4280 25050
rect 4292 24998 4344 25050
rect 4356 24998 4408 25050
rect 4420 24998 4472 25050
rect 34948 24998 35000 25050
rect 35012 24998 35064 25050
rect 35076 24998 35128 25050
rect 35140 24998 35192 25050
rect 2210 24896 2262 24948
rect 2578 24896 2630 24948
rect 7638 24896 7690 24948
rect 7546 24828 7598 24880
rect 8834 24862 8886 24914
rect 9018 24896 9070 24948
rect 21530 24896 21582 24948
rect 23278 24896 23330 24948
rect 23462 24896 23514 24948
rect 45542 24828 45594 24880
rect 45726 24828 45778 24880
rect 2486 24735 2538 24744
rect 2486 24701 2495 24735
rect 2495 24701 2529 24735
rect 2529 24701 2538 24735
rect 2486 24692 2538 24701
rect 20886 24760 20938 24812
rect 8466 24624 8518 24676
rect 8604 24658 8656 24710
rect 20978 24692 21030 24744
rect 9018 24624 9070 24676
rect 21714 24624 21766 24676
rect 19588 24454 19640 24506
rect 19652 24454 19704 24506
rect 19716 24454 19768 24506
rect 19780 24454 19832 24506
rect 50308 24454 50360 24506
rect 50372 24454 50424 24506
rect 50436 24454 50488 24506
rect 50500 24454 50552 24506
rect 8466 24352 8518 24404
rect 21806 24352 21858 24404
rect 2486 24284 2538 24336
rect 28430 24284 28482 24336
rect 43610 24259 43662 24268
rect 43610 24225 43619 24259
rect 43619 24225 43653 24259
rect 43653 24225 43662 24259
rect 43610 24216 43662 24225
rect 7638 24148 7690 24200
rect 32110 24148 32162 24200
rect 56582 24148 56634 24200
rect 56766 24148 56818 24200
rect 12790 24080 12842 24132
rect 20334 24080 20386 24132
rect 6718 24012 6770 24064
rect 4228 23910 4280 23962
rect 4292 23910 4344 23962
rect 4356 23910 4408 23962
rect 4420 23910 4472 23962
rect 34948 23910 35000 23962
rect 35012 23910 35064 23962
rect 35076 23910 35128 23962
rect 35140 23910 35192 23962
rect 7638 23851 7690 23860
rect 7638 23817 7647 23851
rect 7647 23817 7681 23851
rect 7681 23817 7690 23851
rect 7638 23808 7690 23817
rect 8650 23808 8702 23860
rect 8834 23808 8886 23860
rect 12882 23783 12934 23792
rect 12882 23749 12891 23783
rect 12891 23749 12925 23783
rect 12925 23749 12934 23783
rect 12882 23740 12934 23749
rect 27050 23808 27102 23860
rect 13066 23740 13118 23792
rect 8420 23570 8472 23622
rect 12790 23604 12842 23656
rect 18770 23672 18822 23724
rect 20150 23604 20202 23656
rect 8742 23536 8794 23588
rect 12882 23536 12934 23588
rect 32478 23536 32530 23588
rect 20242 23468 20294 23520
rect 19588 23366 19640 23418
rect 19652 23366 19704 23418
rect 19716 23366 19768 23418
rect 19780 23366 19832 23418
rect 50308 23366 50360 23418
rect 50372 23366 50424 23418
rect 50436 23366 50488 23418
rect 50500 23366 50552 23418
rect 26498 22924 26550 22976
rect 26682 22924 26734 22976
rect 4228 22822 4280 22874
rect 4292 22822 4344 22874
rect 4356 22822 4408 22874
rect 4420 22822 4472 22874
rect 34948 22822 35000 22874
rect 35012 22822 35064 22874
rect 35076 22822 35128 22874
rect 35140 22822 35192 22874
rect 18402 22720 18454 22772
rect 33030 22584 33082 22636
rect 18310 22516 18362 22568
rect 25946 22516 25998 22568
rect 18034 22448 18086 22500
rect 18494 22380 18546 22432
rect 19588 22278 19640 22330
rect 19652 22278 19704 22330
rect 19716 22278 19768 22330
rect 19780 22278 19832 22330
rect 50308 22278 50360 22330
rect 50372 22278 50424 22330
rect 50436 22278 50488 22330
rect 50500 22278 50552 22330
rect 33766 22108 33818 22160
rect 13434 21836 13486 21888
rect 50602 21904 50654 21956
rect 35514 21836 35566 21888
rect 47934 21879 47986 21888
rect 47934 21845 47943 21879
rect 47943 21845 47977 21879
rect 47977 21845 47986 21879
rect 47934 21836 47986 21845
rect 4228 21734 4280 21786
rect 4292 21734 4344 21786
rect 4356 21734 4408 21786
rect 4420 21734 4472 21786
rect 34948 21734 35000 21786
rect 35012 21734 35064 21786
rect 35076 21734 35128 21786
rect 35140 21734 35192 21786
rect 17022 21496 17074 21548
rect 16930 21428 16982 21480
rect 42138 21428 42190 21480
rect 8466 21292 8518 21344
rect 8650 21292 8702 21344
rect 16838 21292 16890 21344
rect 19588 21190 19640 21242
rect 19652 21190 19704 21242
rect 19716 21190 19768 21242
rect 19780 21190 19832 21242
rect 50308 21190 50360 21242
rect 50372 21190 50424 21242
rect 50436 21190 50488 21242
rect 50500 21190 50552 21242
rect 18770 20816 18822 20868
rect 19966 20816 20018 20868
rect 4228 20646 4280 20698
rect 4292 20646 4344 20698
rect 4356 20646 4408 20698
rect 4420 20646 4472 20698
rect 34948 20646 35000 20698
rect 35012 20646 35064 20698
rect 35076 20646 35128 20698
rect 35140 20646 35192 20698
rect 8466 20544 8518 20596
rect 48118 20544 48170 20596
rect 9478 20408 9530 20460
rect 10858 20383 10910 20392
rect 8420 20306 8472 20358
rect 10858 20349 10867 20383
rect 10867 20349 10901 20383
rect 10901 20349 10910 20383
rect 10858 20340 10910 20349
rect 48118 20340 48170 20392
rect 16194 20272 16246 20324
rect 14538 20204 14590 20256
rect 19588 20102 19640 20154
rect 19652 20102 19704 20154
rect 19716 20102 19768 20154
rect 19780 20102 19832 20154
rect 50308 20102 50360 20154
rect 50372 20102 50424 20154
rect 50436 20102 50488 20154
rect 50500 20102 50552 20154
rect 8466 20000 8518 20052
rect 16286 20000 16338 20052
rect 5614 19796 5666 19848
rect 10950 19728 11002 19780
rect 27326 19796 27378 19848
rect 49038 19796 49090 19848
rect 26038 19660 26090 19712
rect 27418 19660 27470 19712
rect 4228 19558 4280 19610
rect 4292 19558 4344 19610
rect 4356 19558 4408 19610
rect 4420 19558 4472 19610
rect 34948 19558 35000 19610
rect 35012 19558 35064 19610
rect 35076 19558 35128 19610
rect 35140 19558 35192 19610
rect 5614 19499 5666 19508
rect 5614 19465 5623 19499
rect 5623 19465 5657 19499
rect 5657 19465 5666 19499
rect 5614 19456 5666 19465
rect 8466 19456 8518 19508
rect 21346 19388 21398 19440
rect 26958 19320 27010 19372
rect 37906 19320 37958 19372
rect 37998 19320 38050 19372
rect 51062 19320 51114 19372
rect 51246 19320 51298 19372
rect 7270 19295 7322 19304
rect 7270 19261 7279 19295
rect 7279 19261 7313 19295
rect 7313 19261 7322 19295
rect 7270 19252 7322 19261
rect 8420 19218 8472 19270
rect 21162 19252 21214 19304
rect 27050 19252 27102 19304
rect 20702 19184 20754 19236
rect 23186 19184 23238 19236
rect 8190 19116 8242 19168
rect 8926 19116 8978 19168
rect 13066 19116 13118 19168
rect 19588 19014 19640 19066
rect 19652 19014 19704 19066
rect 19716 19014 19768 19066
rect 19780 19014 19832 19066
rect 50308 19014 50360 19066
rect 50372 19014 50424 19066
rect 50436 19014 50488 19066
rect 50500 19014 50552 19066
rect 8466 18912 8518 18964
rect 10398 18912 10450 18964
rect 8558 18844 8610 18896
rect 16746 18844 16798 18896
rect 27602 18708 27654 18760
rect 27786 18708 27838 18760
rect 7270 18640 7322 18692
rect 17942 18640 17994 18692
rect 2394 18572 2446 18624
rect 47474 18572 47526 18624
rect 4228 18470 4280 18522
rect 4292 18470 4344 18522
rect 4356 18470 4408 18522
rect 4420 18470 4472 18522
rect 34948 18470 35000 18522
rect 35012 18470 35064 18522
rect 35076 18470 35128 18522
rect 35140 18470 35192 18522
rect 7270 18368 7322 18420
rect 8834 18368 8886 18420
rect 9018 18368 9070 18420
rect 14170 18368 14222 18420
rect 13618 18232 13670 18284
rect 11502 18164 11554 18216
rect 51706 18164 51758 18216
rect 33214 18096 33266 18148
rect 40666 18096 40718 18148
rect 44162 18096 44214 18148
rect 12790 18028 12842 18080
rect 19588 17926 19640 17978
rect 19652 17926 19704 17978
rect 19716 17926 19768 17978
rect 19780 17926 19832 17978
rect 50308 17926 50360 17978
rect 50372 17926 50424 17978
rect 50436 17926 50488 17978
rect 50500 17926 50552 17978
rect 27970 17824 28022 17876
rect 8834 17756 8886 17808
rect 56766 17756 56818 17808
rect 8742 17688 8794 17740
rect 55202 17688 55254 17740
rect 1198 17620 1250 17672
rect 27970 17552 28022 17604
rect 39286 17620 39338 17672
rect 19322 17484 19374 17536
rect 24566 17484 24618 17536
rect 38274 17484 38326 17536
rect 48762 17484 48814 17536
rect 4228 17382 4280 17434
rect 4292 17382 4344 17434
rect 4356 17382 4408 17434
rect 4420 17382 4472 17434
rect 34948 17382 35000 17434
rect 35012 17382 35064 17434
rect 35076 17382 35128 17434
rect 35140 17382 35192 17434
rect 8006 17280 8058 17332
rect 8834 17280 8886 17332
rect 7822 17076 7874 17128
rect 9202 17246 9254 17298
rect 23370 17280 23422 17332
rect 33122 17280 33174 17332
rect 8742 17076 8794 17128
rect 24566 17076 24618 17128
rect 24750 17076 24802 17128
rect 19588 16838 19640 16890
rect 19652 16838 19704 16890
rect 19716 16838 19768 16890
rect 19780 16838 19832 16890
rect 50308 16838 50360 16890
rect 50372 16838 50424 16890
rect 50436 16838 50488 16890
rect 50500 16838 50552 16890
rect 8650 16396 8702 16448
rect 51062 16396 51114 16448
rect 4228 16294 4280 16346
rect 4292 16294 4344 16346
rect 4356 16294 4408 16346
rect 4420 16294 4472 16346
rect 34948 16294 35000 16346
rect 35012 16294 35064 16346
rect 35076 16294 35128 16346
rect 35140 16294 35192 16346
rect 8742 16192 8794 16244
rect 36526 16192 36578 16244
rect 8650 16074 8702 16126
rect 24934 16124 24986 16176
rect 24566 16056 24618 16108
rect 3038 15988 3090 16040
rect 15090 15988 15142 16040
rect 34594 16031 34646 16040
rect 34594 15997 34603 16031
rect 34603 15997 34637 16031
rect 34637 15997 34646 16031
rect 34594 15988 34646 15997
rect 34778 15988 34830 16040
rect 24750 15920 24802 15972
rect 24934 15920 24986 15972
rect 8742 15852 8794 15904
rect 15182 15852 15234 15904
rect 19588 15750 19640 15802
rect 19652 15750 19704 15802
rect 19716 15750 19768 15802
rect 19780 15750 19832 15802
rect 50308 15750 50360 15802
rect 50372 15750 50424 15802
rect 50436 15750 50488 15802
rect 50500 15750 50552 15802
rect 50694 15376 50746 15428
rect 45358 15308 45410 15360
rect 45542 15308 45594 15360
rect 48210 15308 48262 15360
rect 4228 15206 4280 15258
rect 4292 15206 4344 15258
rect 4356 15206 4408 15258
rect 4420 15206 4472 15258
rect 34948 15206 35000 15258
rect 35012 15206 35064 15258
rect 35076 15206 35128 15258
rect 35140 15206 35192 15258
rect 8466 15104 8518 15156
rect 8650 15104 8702 15156
rect 35330 15104 35382 15156
rect 13802 15036 13854 15088
rect 18678 15036 18730 15088
rect 8650 14968 8702 15020
rect 48394 14968 48446 15020
rect 2302 14900 2354 14952
rect 8374 14866 8426 14918
rect 29626 14900 29678 14952
rect 46830 14900 46882 14952
rect 19588 14662 19640 14714
rect 19652 14662 19704 14714
rect 19716 14662 19768 14714
rect 19780 14662 19832 14714
rect 50308 14662 50360 14714
rect 50372 14662 50424 14714
rect 50436 14662 50488 14714
rect 50500 14662 50552 14714
rect 18402 14492 18454 14544
rect 18862 14492 18914 14544
rect 44622 14467 44674 14476
rect 44622 14433 44631 14467
rect 44631 14433 44665 14467
rect 44665 14433 44674 14467
rect 44622 14424 44674 14433
rect 6994 14356 7046 14408
rect 25670 14356 25722 14408
rect 7638 14288 7690 14340
rect 25762 14263 25814 14272
rect 25762 14229 25771 14263
rect 25771 14229 25805 14263
rect 25805 14229 25814 14263
rect 25762 14220 25814 14229
rect 45174 14220 45226 14272
rect 52350 14220 52402 14272
rect 4228 14118 4280 14170
rect 4292 14118 4344 14170
rect 4356 14118 4408 14170
rect 4420 14118 4472 14170
rect 34948 14118 35000 14170
rect 35012 14118 35064 14170
rect 35076 14118 35128 14170
rect 35140 14118 35192 14170
rect 6994 14059 7046 14068
rect 6994 14025 7003 14059
rect 7003 14025 7037 14059
rect 7037 14025 7046 14059
rect 6994 14016 7046 14025
rect 10582 14016 10634 14068
rect 25762 14016 25814 14068
rect 40666 13948 40718 14000
rect 32386 13880 32438 13932
rect 8006 13812 8058 13864
rect 12514 13812 12566 13864
rect 45542 13812 45594 13864
rect 49866 13787 49918 13796
rect 49866 13753 49875 13787
rect 49875 13753 49909 13787
rect 49909 13753 49918 13787
rect 49866 13744 49918 13753
rect 19588 13574 19640 13626
rect 19652 13574 19704 13626
rect 19716 13574 19768 13626
rect 19780 13574 19832 13626
rect 50308 13574 50360 13626
rect 50372 13574 50424 13626
rect 50436 13574 50488 13626
rect 50500 13574 50552 13626
rect 3682 13132 3734 13184
rect 17114 13132 17166 13184
rect 4228 13030 4280 13082
rect 4292 13030 4344 13082
rect 4356 13030 4408 13082
rect 4420 13030 4472 13082
rect 34948 13030 35000 13082
rect 35012 13030 35064 13082
rect 35076 13030 35128 13082
rect 35140 13030 35192 13082
rect 8144 12928 8196 12980
rect 17114 12928 17166 12980
rect 44714 12971 44766 12980
rect 44714 12937 44723 12971
rect 44723 12937 44757 12971
rect 44757 12937 44766 12971
rect 44714 12928 44766 12937
rect 21346 12792 21398 12844
rect 21898 12792 21950 12844
rect 10766 12724 10818 12776
rect 23830 12767 23882 12776
rect 23830 12733 23839 12767
rect 23839 12733 23873 12767
rect 23873 12733 23882 12767
rect 23830 12724 23882 12733
rect 21346 12656 21398 12708
rect 42874 12724 42926 12776
rect 51798 12724 51850 12776
rect 19588 12486 19640 12538
rect 19652 12486 19704 12538
rect 19716 12486 19768 12538
rect 19780 12486 19832 12538
rect 50308 12486 50360 12538
rect 50372 12486 50424 12538
rect 50436 12486 50488 12538
rect 50500 12486 50552 12538
rect 21070 12384 21122 12436
rect 11502 12316 11554 12368
rect 13250 12316 13302 12368
rect 7822 12248 7874 12300
rect 26222 12248 26274 12300
rect 48762 12316 48814 12368
rect 49222 12316 49274 12368
rect 6442 12180 6494 12232
rect 6810 12180 6862 12232
rect 6810 12044 6862 12096
rect 26222 12112 26274 12164
rect 40298 12044 40350 12096
rect 44070 12044 44122 12096
rect 4228 11942 4280 11994
rect 4292 11942 4344 11994
rect 4356 11942 4408 11994
rect 4420 11942 4472 11994
rect 34948 11942 35000 11994
rect 35012 11942 35064 11994
rect 35076 11942 35128 11994
rect 35140 11942 35192 11994
rect 11686 11840 11738 11892
rect 15182 11840 15234 11892
rect 6442 11704 6494 11756
rect 6810 11704 6862 11756
rect 8098 11704 8150 11756
rect 26222 11704 26274 11756
rect 37354 11704 37406 11756
rect 19046 11679 19098 11688
rect 19046 11645 19055 11679
rect 19055 11645 19089 11679
rect 19089 11645 19098 11679
rect 19046 11636 19098 11645
rect 24842 11568 24894 11620
rect 26222 11568 26274 11620
rect 37906 11500 37958 11552
rect 59710 11636 59762 11688
rect 58606 11568 58658 11620
rect 19588 11398 19640 11450
rect 19652 11398 19704 11450
rect 19716 11398 19768 11450
rect 19780 11398 19832 11450
rect 50308 11398 50360 11450
rect 50372 11398 50424 11450
rect 50436 11398 50488 11450
rect 50500 11398 50552 11450
rect 9294 10956 9346 11008
rect 33306 10956 33358 11008
rect 4228 10854 4280 10906
rect 4292 10854 4344 10906
rect 4356 10854 4408 10906
rect 4420 10854 4472 10906
rect 34948 10854 35000 10906
rect 35012 10854 35064 10906
rect 35076 10854 35128 10906
rect 35140 10854 35192 10906
rect 24842 10752 24894 10804
rect 26222 10752 26274 10804
rect 29810 10795 29862 10804
rect 29810 10761 29819 10795
rect 29819 10761 29853 10795
rect 29853 10761 29862 10795
rect 29810 10752 29862 10761
rect 9662 10548 9714 10600
rect 9846 10548 9898 10600
rect 26222 10616 26274 10668
rect 38642 10616 38694 10668
rect 24750 10548 24802 10600
rect 9294 10480 9346 10532
rect 19588 10310 19640 10362
rect 19652 10310 19704 10362
rect 19716 10310 19768 10362
rect 19780 10310 19832 10362
rect 50308 10310 50360 10362
rect 50372 10310 50424 10362
rect 50436 10310 50488 10362
rect 50500 10310 50552 10362
rect 9662 10208 9714 10260
rect 34502 10208 34554 10260
rect 21346 10072 21398 10124
rect 24014 10072 24066 10124
rect 2210 10004 2262 10056
rect 10398 9936 10450 9988
rect 10674 9936 10726 9988
rect 24014 9936 24066 9988
rect 3866 9868 3918 9920
rect 21346 9868 21398 9920
rect 32294 9911 32346 9920
rect 32294 9877 32303 9911
rect 32303 9877 32337 9911
rect 32337 9877 32346 9911
rect 32294 9868 32346 9877
rect 50142 9868 50194 9920
rect 4228 9766 4280 9818
rect 4292 9766 4344 9818
rect 4356 9766 4408 9818
rect 4420 9766 4472 9818
rect 34948 9766 35000 9818
rect 35012 9766 35064 9818
rect 35076 9766 35128 9818
rect 35140 9766 35192 9818
rect 6166 9664 6218 9716
rect 17482 9664 17534 9716
rect 32294 9664 32346 9716
rect 41126 9664 41178 9716
rect 44162 9664 44214 9716
rect 6074 9596 6126 9648
rect 7730 9596 7782 9648
rect 8098 9596 8150 9648
rect 10858 9596 10910 9648
rect 11870 9596 11922 9648
rect 7546 9460 7598 9512
rect 7730 9460 7782 9512
rect 8374 9426 8426 9478
rect 10858 9460 10910 9512
rect 11042 9460 11094 9512
rect 31006 9392 31058 9444
rect 19588 9222 19640 9274
rect 19652 9222 19704 9274
rect 19716 9222 19768 9274
rect 19780 9222 19832 9274
rect 50308 9222 50360 9274
rect 50372 9222 50424 9274
rect 50436 9222 50488 9274
rect 50500 9222 50552 9274
rect 8374 9120 8426 9172
rect 29350 9120 29402 9172
rect 2854 8780 2906 8832
rect 48394 8780 48446 8832
rect 4228 8678 4280 8730
rect 4292 8678 4344 8730
rect 4356 8678 4408 8730
rect 4420 8678 4472 8730
rect 34948 8678 35000 8730
rect 35012 8678 35064 8730
rect 35076 8678 35128 8730
rect 35140 8678 35192 8730
rect 24014 8576 24066 8628
rect 26958 8576 27010 8628
rect 28246 8576 28298 8628
rect 48394 8619 48446 8628
rect 48394 8585 48403 8619
rect 48403 8585 48437 8619
rect 48437 8585 48446 8619
rect 48394 8576 48446 8585
rect 3958 8483 4010 8492
rect 3958 8449 3967 8483
rect 3967 8449 4001 8483
rect 4001 8449 4010 8483
rect 3958 8440 4010 8449
rect 8834 8440 8886 8492
rect 26590 8440 26642 8492
rect 26958 8440 27010 8492
rect 40666 8508 40718 8560
rect 41402 8508 41454 8560
rect 8558 8372 8610 8424
rect 20702 8372 20754 8424
rect 21438 8372 21490 8424
rect 10950 8304 11002 8356
rect 40298 8236 40350 8288
rect 47290 8236 47342 8288
rect 19588 8134 19640 8186
rect 19652 8134 19704 8186
rect 19716 8134 19768 8186
rect 19780 8134 19832 8186
rect 50308 8134 50360 8186
rect 50372 8134 50424 8186
rect 50436 8134 50488 8186
rect 50500 8134 50552 8186
rect 21070 8032 21122 8084
rect 21622 8032 21674 8084
rect 22818 7896 22870 7948
rect 23370 7896 23422 7948
rect 15642 7828 15694 7880
rect 16378 7828 16430 7880
rect 22358 7828 22410 7880
rect 22726 7828 22778 7880
rect 12238 7760 12290 7812
rect 15918 7692 15970 7744
rect 16378 7692 16430 7744
rect 21346 7692 21398 7744
rect 21806 7692 21858 7744
rect 22634 7692 22686 7744
rect 22910 7692 22962 7744
rect 25118 7735 25170 7744
rect 25118 7701 25127 7735
rect 25127 7701 25161 7735
rect 25161 7701 25170 7735
rect 25118 7692 25170 7701
rect 25578 7692 25630 7744
rect 25946 7692 25998 7744
rect 46278 7735 46330 7744
rect 46278 7701 46287 7735
rect 46287 7701 46321 7735
rect 46321 7701 46330 7735
rect 46278 7692 46330 7701
rect 4228 7590 4280 7642
rect 4292 7590 4344 7642
rect 4356 7590 4408 7642
rect 4420 7590 4472 7642
rect 34948 7590 35000 7642
rect 35012 7590 35064 7642
rect 35076 7590 35128 7642
rect 35140 7590 35192 7642
rect 15826 7488 15878 7540
rect 16286 7488 16338 7540
rect 18310 7488 18362 7540
rect 18770 7488 18822 7540
rect 19414 7488 19466 7540
rect 20334 7488 20386 7540
rect 23002 7488 23054 7540
rect 23278 7488 23330 7540
rect 28982 7488 29034 7540
rect 29994 7488 30046 7540
rect 31006 7488 31058 7540
rect 46278 7488 46330 7540
rect 25118 7420 25170 7472
rect 34686 7420 34738 7472
rect 8650 7352 8702 7404
rect 23462 7352 23514 7404
rect 8374 7284 8426 7336
rect 16286 7284 16338 7336
rect 24106 7148 24158 7200
rect 19588 7046 19640 7098
rect 19652 7046 19704 7098
rect 19716 7046 19768 7098
rect 19780 7046 19832 7098
rect 50308 7046 50360 7098
rect 50372 7046 50424 7098
rect 50436 7046 50488 7098
rect 50500 7046 50552 7098
rect 8190 6672 8242 6724
rect 10030 6672 10082 6724
rect 5338 6604 5390 6656
rect 8466 6604 8518 6656
rect 10122 6604 10174 6656
rect 4228 6502 4280 6554
rect 4292 6502 4344 6554
rect 4356 6502 4408 6554
rect 4420 6502 4472 6554
rect 34948 6502 35000 6554
rect 35012 6502 35064 6554
rect 35076 6502 35128 6554
rect 35140 6502 35192 6554
rect 8190 6400 8242 6452
rect 8466 6400 8518 6452
rect 17298 6400 17350 6452
rect 18954 6264 19006 6316
rect 10582 6196 10634 6248
rect 26222 6128 26274 6180
rect 14446 6060 14498 6112
rect 19588 5958 19640 6010
rect 19652 5958 19704 6010
rect 19716 5958 19768 6010
rect 19780 5958 19832 6010
rect 50308 5958 50360 6010
rect 50372 5958 50424 6010
rect 50436 5958 50488 6010
rect 50500 5958 50552 6010
rect 1290 5856 1342 5908
rect 8466 5856 8518 5908
rect 20610 5856 20662 5908
rect 4602 5584 4654 5636
rect 14906 5516 14958 5568
rect 4228 5414 4280 5466
rect 4292 5414 4344 5466
rect 4356 5414 4408 5466
rect 4420 5414 4472 5466
rect 34948 5414 35000 5466
rect 35012 5414 35064 5466
rect 35076 5414 35128 5466
rect 35140 5414 35192 5466
rect 8236 5210 8288 5262
rect 12422 5312 12474 5364
rect 11318 5176 11370 5228
rect 8742 5108 8794 5160
rect 15274 5108 15326 5160
rect 8650 4972 8702 5024
rect 20978 4972 21030 5024
rect 21714 4972 21766 5024
rect 19588 4870 19640 4922
rect 19652 4870 19704 4922
rect 19716 4870 19768 4922
rect 19780 4870 19832 4922
rect 50308 4870 50360 4922
rect 50372 4870 50424 4922
rect 50436 4870 50488 4922
rect 50500 4870 50552 4922
rect 12790 4768 12842 4820
rect 12974 4768 13026 4820
rect 17022 4768 17074 4820
rect 17390 4768 17442 4820
rect 40206 4768 40258 4820
rect 41126 4768 41178 4820
rect 30086 4632 30138 4684
rect 37262 4632 37314 4684
rect 23830 4496 23882 4548
rect 31650 4496 31702 4548
rect 38274 4496 38326 4548
rect 47014 4496 47066 4548
rect 7454 4428 7506 4480
rect 31834 4428 31886 4480
rect 41034 4428 41086 4480
rect 4228 4326 4280 4378
rect 4292 4326 4344 4378
rect 4356 4326 4408 4378
rect 4420 4326 4472 4378
rect 34948 4326 35000 4378
rect 35012 4326 35064 4378
rect 35076 4326 35128 4378
rect 35140 4326 35192 4378
rect 7454 4267 7506 4276
rect 7454 4233 7463 4267
rect 7463 4233 7497 4267
rect 7497 4233 7506 4267
rect 7454 4224 7506 4233
rect 9110 4224 9162 4276
rect 21162 4224 21214 4276
rect 22266 4224 22318 4276
rect 25026 4224 25078 4276
rect 18954 4156 19006 4208
rect 27418 4156 27470 4208
rect 3682 4088 3734 4140
rect 3958 4088 4010 4140
rect 4694 4088 4746 4140
rect 5154 4088 5206 4140
rect 6166 4088 6218 4140
rect 6718 4088 6770 4140
rect 7638 4088 7690 4140
rect 8006 4088 8058 4140
rect 8098 4088 8150 4140
rect 9846 4088 9898 4140
rect 10766 4088 10818 4140
rect 11686 4088 11738 4140
rect 12330 4088 12382 4140
rect 13066 4088 13118 4140
rect 13342 4088 13394 4140
rect 13434 4088 13486 4140
rect 13710 4088 13762 4140
rect 14538 4088 14590 4140
rect 15458 4088 15510 4140
rect 16010 4088 16062 4140
rect 16470 4088 16522 4140
rect 17114 4088 17166 4140
rect 17850 4088 17902 4140
rect 18862 4088 18914 4140
rect 19322 4088 19374 4140
rect 20058 4088 20110 4140
rect 20426 4088 20478 4140
rect 21254 4088 21306 4140
rect 22634 4088 22686 4140
rect 24290 4088 24342 4140
rect 25026 4088 25078 4140
rect 25210 4088 25262 4140
rect 26130 4088 26182 4140
rect 26314 4088 26366 4140
rect 27510 4088 27562 4140
rect 28522 4088 28574 4140
rect 29626 4088 29678 4140
rect 3222 4020 3274 4072
rect 4050 4020 4102 4072
rect 5062 4020 5114 4072
rect 5430 4020 5482 4072
rect 11318 4020 11370 4072
rect 12054 4020 12106 4072
rect 13802 4020 13854 4072
rect 14998 4020 15050 4072
rect 19966 4020 20018 4072
rect 20794 4020 20846 4072
rect 22818 4020 22870 4072
rect 24842 4020 24894 4072
rect 27050 4020 27102 4072
rect 4970 3952 5022 4004
rect 6902 3952 6954 4004
rect 6258 3884 6310 3936
rect 12790 3952 12842 4004
rect 13526 3952 13578 4004
rect 16838 3952 16890 4004
rect 17850 3952 17902 4004
rect 20150 3952 20202 4004
rect 21162 3952 21214 4004
rect 21254 3952 21306 4004
rect 22542 3952 22594 4004
rect 25486 3952 25538 4004
rect 28154 3952 28206 4004
rect 28890 4020 28942 4072
rect 30178 4020 30230 4072
rect 31650 4088 31702 4140
rect 43150 4224 43202 4276
rect 32846 3952 32898 4004
rect 33950 4020 34002 4072
rect 34410 4020 34462 4072
rect 34594 4020 34646 4072
rect 37998 4020 38050 4072
rect 38550 4020 38602 4072
rect 39654 4156 39706 4208
rect 39746 4020 39798 4072
rect 46738 4088 46790 4140
rect 50786 4088 50838 4140
rect 51798 4088 51850 4140
rect 54190 4088 54242 4140
rect 10674 3884 10726 3936
rect 14446 3884 14498 3936
rect 15734 3884 15786 3936
rect 31742 3884 31794 3936
rect 31834 3884 31886 3936
rect 33214 3884 33266 3936
rect 35238 3884 35290 3936
rect 36526 3884 36578 3936
rect 36618 3884 36670 3936
rect 39102 3884 39154 3936
rect 39194 3884 39246 3936
rect 40574 3884 40626 3936
rect 40758 3884 40810 3936
rect 51614 4020 51666 4072
rect 49774 3952 49826 4004
rect 50970 3952 51022 4004
rect 48946 3884 48998 3936
rect 56766 3884 56818 3936
rect 19588 3782 19640 3834
rect 19652 3782 19704 3834
rect 19716 3782 19768 3834
rect 19780 3782 19832 3834
rect 50308 3782 50360 3834
rect 50372 3782 50424 3834
rect 50436 3782 50488 3834
rect 50500 3782 50552 3834
rect 8374 3680 8426 3732
rect 11778 3680 11830 3732
rect 11870 3680 11922 3732
rect 7270 3612 7322 3664
rect 11042 3612 11094 3664
rect 12882 3612 12934 3664
rect 14814 3612 14866 3664
rect 23186 3680 23238 3732
rect 24290 3680 24342 3732
rect 27510 3680 27562 3732
rect 28982 3680 29034 3732
rect 31742 3680 31794 3732
rect 32938 3680 32990 3732
rect 33030 3680 33082 3732
rect 39194 3680 39246 3732
rect 31834 3612 31886 3664
rect 186 3544 238 3596
rect 1014 3544 1066 3596
rect 1382 3544 1434 3596
rect 2394 3544 2446 3596
rect 6350 3544 6402 3596
rect 14354 3544 14406 3596
rect 17298 3544 17350 3596
rect 40390 3612 40442 3664
rect 36618 3544 36670 3596
rect 38642 3544 38694 3596
rect 38734 3544 38786 3596
rect 39930 3544 39982 3596
rect 5338 3476 5390 3528
rect 31650 3476 31702 3528
rect 3038 3408 3090 3460
rect 37814 3476 37866 3528
rect 48670 3680 48722 3732
rect 49038 3680 49090 3732
rect 42046 3612 42098 3664
rect 46922 3612 46974 3664
rect 47474 3612 47526 3664
rect 49958 3612 50010 3664
rect 47934 3544 47986 3596
rect 51246 3612 51298 3664
rect 51706 3680 51758 3732
rect 59342 3680 59394 3732
rect 57502 3612 57554 3664
rect 50142 3544 50194 3596
rect 54926 3544 54978 3596
rect 47290 3476 47342 3528
rect 48302 3476 48354 3528
rect 39930 3408 39982 3460
rect 45726 3408 45778 3460
rect 46830 3408 46882 3460
rect 47014 3408 47066 3460
rect 53822 3476 53874 3528
rect 14630 3340 14682 3392
rect 21254 3340 21306 3392
rect 21438 3340 21490 3392
rect 22082 3340 22134 3392
rect 23094 3340 23146 3392
rect 23922 3340 23974 3392
rect 24382 3340 24434 3392
rect 27050 3340 27102 3392
rect 28338 3340 28390 3392
rect 31098 3340 31150 3392
rect 31650 3340 31702 3392
rect 34594 3340 34646 3392
rect 36526 3340 36578 3392
rect 46094 3340 46146 3392
rect 47566 3340 47618 3392
rect 55294 3340 55346 3392
rect 4228 3238 4280 3290
rect 4292 3238 4344 3290
rect 4356 3238 4408 3290
rect 4420 3238 4472 3290
rect 34948 3238 35000 3290
rect 35012 3238 35064 3290
rect 35076 3238 35128 3290
rect 35140 3238 35192 3290
rect 6074 3136 6126 3188
rect 10858 3136 10910 3188
rect 17298 3136 17350 3188
rect 18586 3179 18638 3188
rect 18586 3145 18595 3179
rect 18595 3145 18629 3179
rect 18629 3145 18638 3179
rect 18586 3136 18638 3145
rect 22542 3136 22594 3188
rect 36158 3136 36210 3188
rect 38366 3136 38418 3188
rect 41034 3136 41086 3188
rect 41310 3136 41362 3188
rect 45266 3136 45318 3188
rect 46922 3136 46974 3188
rect 50142 3136 50194 3188
rect 50602 3136 50654 3188
rect 58974 3136 59026 3188
rect 8834 3068 8886 3120
rect 19046 3068 19098 3120
rect 23370 3068 23422 3120
rect 25946 3068 25998 3120
rect 26958 3068 27010 3120
rect 29626 3068 29678 3120
rect 38090 3068 38142 3120
rect 47934 3068 47986 3120
rect 49682 3068 49734 3120
rect 50510 3068 50562 3120
rect 50694 3068 50746 3120
rect 58238 3068 58290 3120
rect 2670 3000 2722 3052
rect 8466 3000 8518 3052
rect 16286 3000 16338 3052
rect 18586 3000 18638 3052
rect 21070 3000 21122 3052
rect 23738 3000 23790 3052
rect 24198 3000 24250 3052
rect 27418 3000 27470 3052
rect 27878 3000 27930 3052
rect 28338 3000 28390 3052
rect 29534 3000 29586 3052
rect 36526 3000 36578 3052
rect 38182 3000 38234 3052
rect 20702 2932 20754 2984
rect 23370 2932 23422 2984
rect 26222 2932 26274 2984
rect 29350 2932 29402 2984
rect 29442 2932 29494 2984
rect 39470 2932 39522 2984
rect 39746 3000 39798 3052
rect 41218 3000 41270 3052
rect 41402 3000 41454 3052
rect 51982 3000 52034 3052
rect 54558 3000 54610 3052
rect 55110 3000 55162 3052
rect 42782 2932 42834 2984
rect 45266 2932 45318 2984
rect 49038 2932 49090 2984
rect 22358 2864 22410 2916
rect 26682 2864 26734 2916
rect 28430 2864 28482 2916
rect 9570 2796 9622 2848
rect 12054 2796 12106 2848
rect 27142 2796 27194 2848
rect 30822 2796 30874 2848
rect 31098 2864 31150 2916
rect 33582 2864 33634 2916
rect 33674 2864 33726 2916
rect 34318 2796 34370 2848
rect 34594 2864 34646 2916
rect 39838 2864 39890 2916
rect 41310 2864 41362 2916
rect 41678 2864 41730 2916
rect 42138 2864 42190 2916
rect 40758 2796 40810 2848
rect 40850 2796 40902 2848
rect 44254 2796 44306 2848
rect 44806 2864 44858 2916
rect 56398 2932 56450 2984
rect 50786 2864 50838 2916
rect 53454 2864 53506 2916
rect 49682 2796 49734 2848
rect 50050 2796 50102 2848
rect 57870 2796 57922 2848
rect 19588 2694 19640 2746
rect 19652 2694 19704 2746
rect 19716 2694 19768 2746
rect 19780 2694 19832 2746
rect 50308 2694 50360 2746
rect 50372 2694 50424 2746
rect 50436 2694 50488 2746
rect 50500 2694 50552 2746
rect 22450 2592 22502 2644
rect 22818 2592 22870 2644
rect 22910 2592 22962 2644
rect 23186 2592 23238 2644
rect 25670 2592 25722 2644
rect 27786 2592 27838 2644
rect 30822 2592 30874 2644
rect 32478 2592 32530 2644
rect 39930 2592 39982 2644
rect 40850 2592 40902 2644
rect 40390 2524 40442 2576
rect 42414 2524 42466 2576
rect 48486 2524 48538 2576
rect 53086 2524 53138 2576
rect 9570 2456 9622 2508
rect 12422 2456 12474 2508
rect 13158 2456 13210 2508
rect 50050 2320 50102 2372
rect 14538 2252 14590 2304
rect 4228 2150 4280 2202
rect 4292 2150 4344 2202
rect 4356 2150 4408 2202
rect 4420 2150 4472 2202
rect 34948 2150 35000 2202
rect 35012 2150 35064 2202
rect 35076 2150 35128 2202
rect 35140 2150 35192 2202
rect 30638 2048 30690 2100
rect 31282 2048 31334 2100
rect 30178 1980 30230 2032
rect 36526 1980 36578 2032
rect 29074 1844 29126 1896
rect 35790 1844 35842 1896
rect 39838 1708 39890 1760
rect 41310 1708 41362 1760
rect 38826 1572 38878 1624
rect 39838 1572 39890 1624
rect 17942 1368 17994 1420
rect 18218 1368 18270 1420
rect 19690 1368 19742 1420
rect 20518 1368 20570 1420
rect 29350 1368 29402 1420
rect 30270 1368 30322 1420
rect 49958 1368 50010 1420
rect 50878 1368 50930 1420
rect 29166 892 29218 944
rect 29258 892 29310 944
<< metal2 >>
rect 184 59200 240 60000
rect 644 59200 700 60000
rect 1196 59200 1252 60000
rect 1748 59200 1804 60000
rect 2208 59200 2264 60000
rect 2760 59200 2816 60000
rect 3312 59200 3368 60000
rect 3864 59200 3920 60000
rect 4324 59200 4380 60000
rect 4876 59200 4932 60000
rect 5428 59200 5484 60000
rect 5888 59200 5944 60000
rect 6440 59200 6496 60000
rect 6992 59200 7048 60000
rect 7544 59200 7600 60000
rect 8004 59200 8060 60000
rect 8556 59200 8612 60000
rect 9108 59200 9164 60000
rect 9568 59200 9624 60000
rect 10120 59200 10176 60000
rect 10672 59200 10728 60000
rect 11224 59200 11280 60000
rect 11684 59200 11740 60000
rect 12236 59200 12292 60000
rect 12788 59200 12844 60000
rect 13248 59200 13304 60000
rect 13800 59200 13856 60000
rect 14352 59200 14408 60000
rect 14904 59200 14960 60000
rect 15364 59200 15420 60000
rect 15916 59200 15972 60000
rect 16468 59200 16524 60000
rect 17020 59200 17076 60000
rect 17480 59200 17536 60000
rect 18032 59200 18088 60000
rect 18584 59200 18640 60000
rect 19044 59200 19100 60000
rect 19596 59200 19652 60000
rect 20148 59200 20204 60000
rect 20700 59200 20756 60000
rect 21160 59200 21216 60000
rect 21712 59200 21768 60000
rect 22264 59200 22320 60000
rect 22724 59200 22780 60000
rect 23276 59200 23332 60000
rect 23828 59200 23884 60000
rect 24380 59200 24436 60000
rect 24840 59200 24896 60000
rect 25392 59200 25448 60000
rect 25944 59200 26000 60000
rect 26404 59200 26460 60000
rect 26956 59200 27012 60000
rect 27508 59200 27564 60000
rect 28060 59200 28116 60000
rect 28520 59200 28576 60000
rect 29072 59200 29128 60000
rect 29624 59200 29680 60000
rect 30176 59200 30232 60000
rect 30636 59200 30692 60000
rect 31188 59200 31244 60000
rect 31740 59200 31796 60000
rect 32200 59200 32256 60000
rect 32752 59200 32808 60000
rect 33304 59200 33360 60000
rect 33856 59200 33912 60000
rect 34316 59200 34372 60000
rect 34868 59200 34924 60000
rect 35420 59200 35476 60000
rect 35880 59200 35936 60000
rect 36432 59200 36488 60000
rect 36984 59200 37040 60000
rect 37536 59200 37592 60000
rect 37996 59200 38052 60000
rect 38548 59200 38604 60000
rect 39100 59200 39156 60000
rect 39560 59200 39616 60000
rect 40112 59200 40168 60000
rect 40664 59200 40720 60000
rect 41216 59200 41272 60000
rect 41676 59200 41732 60000
rect 42228 59200 42284 60000
rect 42780 59200 42836 60000
rect 43240 59200 43296 60000
rect 43792 59200 43848 60000
rect 44344 59200 44400 60000
rect 44896 59200 44952 60000
rect 45356 59200 45412 60000
rect 45908 59200 45964 60000
rect 46460 59200 46516 60000
rect 47012 59200 47068 60000
rect 47472 59200 47528 60000
rect 48024 59200 48080 60000
rect 48576 59200 48632 60000
rect 49036 59200 49092 60000
rect 49588 59200 49644 60000
rect 50140 59200 50196 60000
rect 50692 59200 50748 60000
rect 51152 59200 51208 60000
rect 51704 59200 51760 60000
rect 52256 59200 52312 60000
rect 52716 59200 52772 60000
rect 53268 59200 53324 60000
rect 53820 59200 53876 60000
rect 54372 59200 54428 60000
rect 54832 59200 54888 60000
rect 55384 59200 55440 60000
rect 55936 59200 55992 60000
rect 56396 59200 56452 60000
rect 56948 59200 57004 60000
rect 57500 59200 57556 60000
rect 58052 59200 58108 60000
rect 58512 59200 58568 60000
rect 59064 59200 59120 60000
rect 59616 59200 59672 60000
rect 198 56438 226 59200
rect 658 56506 686 59200
rect 1210 57202 1238 59200
rect 1118 57174 1238 57202
rect 646 56500 698 56506
rect 646 56442 698 56448
rect 186 56432 238 56438
rect 186 56374 238 56380
rect 1118 37126 1146 57174
rect 1762 56506 1790 59200
rect 2222 59106 2250 59200
rect 2222 59078 2618 59106
rect 1198 56500 1250 56506
rect 1198 56442 1250 56448
rect 1750 56500 1802 56506
rect 1750 56442 1802 56448
rect 1106 37120 1158 37126
rect 1106 37062 1158 37068
rect 1106 34944 1158 34950
rect 1106 34886 1158 34892
rect 1014 29776 1066 29782
rect 1014 29718 1066 29724
rect 1026 3602 1054 29718
rect 186 3596 238 3602
rect 186 3538 238 3544
rect 1014 3596 1066 3602
rect 1014 3538 1066 3544
rect 198 800 226 3538
rect 1118 3482 1146 34886
rect 1210 17678 1238 56442
rect 1290 56432 1342 56438
rect 1290 56374 1342 56380
rect 1198 17672 1250 17678
rect 1198 17614 1250 17620
rect 1302 5914 1330 56374
rect 2486 32564 2538 32570
rect 2486 32506 2538 32512
rect 2210 24948 2262 24954
rect 2210 24890 2262 24896
rect 2222 10062 2250 24890
rect 2498 24834 2526 32506
rect 2590 24954 2618 59078
rect 2670 56500 2722 56506
rect 2670 56442 2722 56448
rect 2578 24948 2630 24954
rect 2578 24890 2630 24896
rect 2498 24806 2618 24834
rect 2486 24744 2538 24750
rect 2486 24686 2538 24692
rect 2498 24342 2526 24686
rect 2486 24336 2538 24342
rect 2486 24278 2538 24284
rect 2590 21434 2618 24806
rect 2498 21406 2618 21434
rect 2394 18624 2446 18630
rect 2394 18566 2446 18572
rect 2302 14952 2354 14958
rect 2302 14894 2354 14900
rect 2210 10056 2262 10062
rect 2210 9998 2262 10004
rect 1290 5908 1342 5914
rect 1290 5850 1342 5856
rect 1382 3596 1434 3602
rect 1382 3538 1434 3544
rect 934 3454 1146 3482
rect 934 800 962 3454
rect 1394 800 1422 3538
rect 2314 898 2342 14894
rect 2406 3602 2434 18566
rect 2394 3596 2446 3602
rect 2394 3538 2446 3544
rect 2498 3482 2526 21406
rect 1946 870 2342 898
rect 2406 3454 2526 3482
rect 1946 800 1974 870
rect 2406 800 2434 3454
rect 2682 3058 2710 56442
rect 2774 55282 2802 59200
rect 2762 55276 2814 55282
rect 2762 55218 2814 55224
rect 3878 55162 3906 59200
rect 4338 59158 4366 59200
rect 4326 59152 4378 59158
rect 4326 59094 4378 59100
rect 4202 57692 4498 57712
rect 4258 57690 4282 57692
rect 4338 57690 4362 57692
rect 4418 57690 4442 57692
rect 4280 57638 4282 57690
rect 4344 57638 4356 57690
rect 4418 57638 4420 57690
rect 4258 57636 4282 57638
rect 4338 57636 4362 57638
rect 4418 57636 4442 57638
rect 4202 57616 4498 57636
rect 4202 56604 4498 56624
rect 4258 56602 4282 56604
rect 4338 56602 4362 56604
rect 4418 56602 4442 56604
rect 4280 56550 4282 56602
rect 4344 56550 4356 56602
rect 4418 56550 4420 56602
rect 4258 56548 4282 56550
rect 4338 56548 4362 56550
rect 4418 56548 4442 56550
rect 4202 56528 4498 56548
rect 4050 56228 4102 56234
rect 4050 56170 4102 56176
rect 3958 55276 4010 55282
rect 3958 55218 4010 55224
rect 3694 55134 3906 55162
rect 3694 28422 3722 55134
rect 3970 55026 3998 55218
rect 3878 54998 3998 55026
rect 3774 36712 3826 36718
rect 3774 36654 3826 36660
rect 3682 28416 3734 28422
rect 3682 28358 3734 28364
rect 3038 16040 3090 16046
rect 3038 15982 3090 15988
rect 2854 8832 2906 8838
rect 2854 8774 2906 8780
rect 2670 3052 2722 3058
rect 2670 2994 2722 3000
rect 2866 800 2894 8774
rect 3050 3466 3078 15982
rect 3682 13184 3734 13190
rect 3682 13126 3734 13132
rect 3694 4146 3722 13126
rect 3682 4140 3734 4146
rect 3682 4082 3734 4088
rect 3222 4072 3274 4078
rect 3222 4014 3274 4020
rect 3038 3460 3090 3466
rect 3038 3402 3090 3408
rect 3234 800 3262 4014
rect 3786 2666 3814 36654
rect 3878 9926 3906 54998
rect 4062 54754 4090 56170
rect 4202 55516 4498 55536
rect 4258 55514 4282 55516
rect 4338 55514 4362 55516
rect 4418 55514 4442 55516
rect 4280 55462 4282 55514
rect 4344 55462 4356 55514
rect 4418 55462 4420 55514
rect 4258 55460 4282 55462
rect 4338 55460 4362 55462
rect 4418 55460 4442 55462
rect 4202 55440 4498 55460
rect 4890 55350 4918 59200
rect 4878 55344 4930 55350
rect 4878 55286 4930 55292
rect 3970 54726 4090 54754
rect 3866 9920 3918 9926
rect 3866 9862 3918 9868
rect 3970 8498 3998 54726
rect 4050 54528 4102 54534
rect 4050 54470 4102 54476
rect 3958 8492 4010 8498
rect 3958 8434 4010 8440
rect 3958 4140 4010 4146
rect 3958 4082 4010 4088
rect 3602 2638 3814 2666
rect 3602 800 3630 2638
rect 3970 800 3998 4082
rect 4062 4078 4090 54470
rect 4202 54428 4498 54448
rect 4258 54426 4282 54428
rect 4338 54426 4362 54428
rect 4418 54426 4442 54428
rect 4280 54374 4282 54426
rect 4344 54374 4356 54426
rect 4418 54374 4420 54426
rect 4258 54372 4282 54374
rect 4338 54372 4362 54374
rect 4418 54372 4442 54374
rect 4202 54352 4498 54372
rect 4202 53340 4498 53360
rect 4258 53338 4282 53340
rect 4338 53338 4362 53340
rect 4418 53338 4442 53340
rect 4280 53286 4282 53338
rect 4344 53286 4356 53338
rect 4418 53286 4420 53338
rect 4258 53284 4282 53286
rect 4338 53284 4362 53286
rect 4418 53284 4442 53286
rect 4202 53264 4498 53284
rect 5062 52420 5114 52426
rect 5062 52362 5114 52368
rect 4202 52252 4498 52272
rect 4258 52250 4282 52252
rect 4338 52250 4362 52252
rect 4418 52250 4442 52252
rect 4280 52198 4282 52250
rect 4344 52198 4356 52250
rect 4418 52198 4420 52250
rect 4258 52196 4282 52198
rect 4338 52196 4362 52198
rect 4418 52196 4442 52198
rect 4202 52176 4498 52196
rect 4202 51164 4498 51184
rect 4258 51162 4282 51164
rect 4338 51162 4362 51164
rect 4418 51162 4442 51164
rect 4280 51110 4282 51162
rect 4344 51110 4356 51162
rect 4418 51110 4420 51162
rect 4258 51108 4282 51110
rect 4338 51108 4362 51110
rect 4418 51108 4442 51110
rect 4202 51088 4498 51108
rect 4202 50076 4498 50096
rect 4258 50074 4282 50076
rect 4338 50074 4362 50076
rect 4418 50074 4442 50076
rect 4280 50022 4282 50074
rect 4344 50022 4356 50074
rect 4418 50022 4420 50074
rect 4258 50020 4282 50022
rect 4338 50020 4362 50022
rect 4418 50020 4442 50022
rect 4202 50000 4498 50020
rect 4202 48988 4498 49008
rect 4258 48986 4282 48988
rect 4338 48986 4362 48988
rect 4418 48986 4442 48988
rect 4280 48934 4282 48986
rect 4344 48934 4356 48986
rect 4418 48934 4420 48986
rect 4258 48932 4282 48934
rect 4338 48932 4362 48934
rect 4418 48932 4442 48934
rect 4202 48912 4498 48932
rect 4202 47900 4498 47920
rect 4258 47898 4282 47900
rect 4338 47898 4362 47900
rect 4418 47898 4442 47900
rect 4280 47846 4282 47898
rect 4344 47846 4356 47898
rect 4418 47846 4420 47898
rect 4258 47844 4282 47846
rect 4338 47844 4362 47846
rect 4418 47844 4442 47846
rect 4202 47824 4498 47844
rect 4202 46812 4498 46832
rect 4258 46810 4282 46812
rect 4338 46810 4362 46812
rect 4418 46810 4442 46812
rect 4280 46758 4282 46810
rect 4344 46758 4356 46810
rect 4418 46758 4420 46810
rect 4258 46756 4282 46758
rect 4338 46756 4362 46758
rect 4418 46756 4442 46758
rect 4202 46736 4498 46756
rect 4202 45724 4498 45744
rect 4258 45722 4282 45724
rect 4338 45722 4362 45724
rect 4418 45722 4442 45724
rect 4280 45670 4282 45722
rect 4344 45670 4356 45722
rect 4418 45670 4420 45722
rect 4258 45668 4282 45670
rect 4338 45668 4362 45670
rect 4418 45668 4442 45670
rect 4202 45648 4498 45668
rect 4202 44636 4498 44656
rect 4258 44634 4282 44636
rect 4338 44634 4362 44636
rect 4418 44634 4442 44636
rect 4280 44582 4282 44634
rect 4344 44582 4356 44634
rect 4418 44582 4420 44634
rect 4258 44580 4282 44582
rect 4338 44580 4362 44582
rect 4418 44580 4442 44582
rect 4202 44560 4498 44580
rect 4202 43548 4498 43568
rect 4258 43546 4282 43548
rect 4338 43546 4362 43548
rect 4418 43546 4442 43548
rect 4280 43494 4282 43546
rect 4344 43494 4356 43546
rect 4418 43494 4420 43546
rect 4258 43492 4282 43494
rect 4338 43492 4362 43494
rect 4418 43492 4442 43494
rect 4202 43472 4498 43492
rect 4202 42460 4498 42480
rect 4258 42458 4282 42460
rect 4338 42458 4362 42460
rect 4418 42458 4442 42460
rect 4280 42406 4282 42458
rect 4344 42406 4356 42458
rect 4418 42406 4420 42458
rect 4258 42404 4282 42406
rect 4338 42404 4362 42406
rect 4418 42404 4442 42406
rect 4202 42384 4498 42404
rect 4202 41372 4498 41392
rect 4258 41370 4282 41372
rect 4338 41370 4362 41372
rect 4418 41370 4442 41372
rect 4280 41318 4282 41370
rect 4344 41318 4356 41370
rect 4418 41318 4420 41370
rect 4258 41316 4282 41318
rect 4338 41316 4362 41318
rect 4418 41316 4442 41318
rect 4202 41296 4498 41316
rect 4202 40284 4498 40304
rect 4258 40282 4282 40284
rect 4338 40282 4362 40284
rect 4418 40282 4442 40284
rect 4280 40230 4282 40282
rect 4344 40230 4356 40282
rect 4418 40230 4420 40282
rect 4258 40228 4282 40230
rect 4338 40228 4362 40230
rect 4418 40228 4442 40230
rect 4202 40208 4498 40228
rect 4970 40112 5022 40118
rect 4970 40054 5022 40060
rect 4202 39196 4498 39216
rect 4258 39194 4282 39196
rect 4338 39194 4362 39196
rect 4418 39194 4442 39196
rect 4280 39142 4282 39194
rect 4344 39142 4356 39194
rect 4418 39142 4420 39194
rect 4258 39140 4282 39142
rect 4338 39140 4362 39142
rect 4418 39140 4442 39142
rect 4202 39120 4498 39140
rect 4202 38108 4498 38128
rect 4258 38106 4282 38108
rect 4338 38106 4362 38108
rect 4418 38106 4442 38108
rect 4280 38054 4282 38106
rect 4344 38054 4356 38106
rect 4418 38054 4420 38106
rect 4258 38052 4282 38054
rect 4338 38052 4362 38054
rect 4418 38052 4442 38054
rect 4202 38032 4498 38052
rect 4202 37020 4498 37040
rect 4258 37018 4282 37020
rect 4338 37018 4362 37020
rect 4418 37018 4442 37020
rect 4280 36966 4282 37018
rect 4344 36966 4356 37018
rect 4418 36966 4420 37018
rect 4258 36964 4282 36966
rect 4338 36964 4362 36966
rect 4418 36964 4442 36966
rect 4202 36944 4498 36964
rect 4202 35932 4498 35952
rect 4258 35930 4282 35932
rect 4338 35930 4362 35932
rect 4418 35930 4442 35932
rect 4280 35878 4282 35930
rect 4344 35878 4356 35930
rect 4418 35878 4420 35930
rect 4258 35876 4282 35878
rect 4338 35876 4362 35878
rect 4418 35876 4442 35878
rect 4202 35856 4498 35876
rect 4202 34844 4498 34864
rect 4258 34842 4282 34844
rect 4338 34842 4362 34844
rect 4418 34842 4442 34844
rect 4280 34790 4282 34842
rect 4344 34790 4356 34842
rect 4418 34790 4420 34842
rect 4258 34788 4282 34790
rect 4338 34788 4362 34790
rect 4418 34788 4442 34790
rect 4202 34768 4498 34788
rect 4202 33756 4498 33776
rect 4258 33754 4282 33756
rect 4338 33754 4362 33756
rect 4418 33754 4442 33756
rect 4280 33702 4282 33754
rect 4344 33702 4356 33754
rect 4418 33702 4420 33754
rect 4258 33700 4282 33702
rect 4338 33700 4362 33702
rect 4418 33700 4442 33702
rect 4202 33680 4498 33700
rect 4202 32668 4498 32688
rect 4258 32666 4282 32668
rect 4338 32666 4362 32668
rect 4418 32666 4442 32668
rect 4280 32614 4282 32666
rect 4344 32614 4356 32666
rect 4418 32614 4420 32666
rect 4258 32612 4282 32614
rect 4338 32612 4362 32614
rect 4418 32612 4442 32614
rect 4202 32592 4498 32612
rect 4202 31580 4498 31600
rect 4258 31578 4282 31580
rect 4338 31578 4362 31580
rect 4418 31578 4442 31580
rect 4280 31526 4282 31578
rect 4344 31526 4356 31578
rect 4418 31526 4420 31578
rect 4258 31524 4282 31526
rect 4338 31524 4362 31526
rect 4418 31524 4442 31526
rect 4202 31504 4498 31524
rect 4202 30492 4498 30512
rect 4258 30490 4282 30492
rect 4338 30490 4362 30492
rect 4418 30490 4442 30492
rect 4280 30438 4282 30490
rect 4344 30438 4356 30490
rect 4418 30438 4420 30490
rect 4258 30436 4282 30438
rect 4338 30436 4362 30438
rect 4418 30436 4442 30438
rect 4202 30416 4498 30436
rect 4202 29404 4498 29424
rect 4258 29402 4282 29404
rect 4338 29402 4362 29404
rect 4418 29402 4442 29404
rect 4280 29350 4282 29402
rect 4344 29350 4356 29402
rect 4418 29350 4420 29402
rect 4258 29348 4282 29350
rect 4338 29348 4362 29350
rect 4418 29348 4442 29350
rect 4202 29328 4498 29348
rect 4202 28316 4498 28336
rect 4258 28314 4282 28316
rect 4338 28314 4362 28316
rect 4418 28314 4442 28316
rect 4280 28262 4282 28314
rect 4344 28262 4356 28314
rect 4418 28262 4420 28314
rect 4258 28260 4282 28262
rect 4338 28260 4362 28262
rect 4418 28260 4442 28262
rect 4202 28240 4498 28260
rect 4202 27228 4498 27248
rect 4258 27226 4282 27228
rect 4338 27226 4362 27228
rect 4418 27226 4442 27228
rect 4280 27174 4282 27226
rect 4344 27174 4356 27226
rect 4418 27174 4420 27226
rect 4258 27172 4282 27174
rect 4338 27172 4362 27174
rect 4418 27172 4442 27174
rect 4202 27152 4498 27172
rect 4202 26140 4498 26160
rect 4258 26138 4282 26140
rect 4338 26138 4362 26140
rect 4418 26138 4442 26140
rect 4280 26086 4282 26138
rect 4344 26086 4356 26138
rect 4418 26086 4420 26138
rect 4258 26084 4282 26086
rect 4338 26084 4362 26086
rect 4418 26084 4442 26086
rect 4202 26064 4498 26084
rect 4202 25052 4498 25072
rect 4258 25050 4282 25052
rect 4338 25050 4362 25052
rect 4418 25050 4442 25052
rect 4280 24998 4282 25050
rect 4344 24998 4356 25050
rect 4418 24998 4420 25050
rect 4258 24996 4282 24998
rect 4338 24996 4362 24998
rect 4418 24996 4442 24998
rect 4202 24976 4498 24996
rect 4202 23964 4498 23984
rect 4258 23962 4282 23964
rect 4338 23962 4362 23964
rect 4418 23962 4442 23964
rect 4280 23910 4282 23962
rect 4344 23910 4356 23962
rect 4418 23910 4420 23962
rect 4258 23908 4282 23910
rect 4338 23908 4362 23910
rect 4418 23908 4442 23910
rect 4202 23888 4498 23908
rect 4202 22876 4498 22896
rect 4258 22874 4282 22876
rect 4338 22874 4362 22876
rect 4418 22874 4442 22876
rect 4280 22822 4282 22874
rect 4344 22822 4356 22874
rect 4418 22822 4420 22874
rect 4258 22820 4282 22822
rect 4338 22820 4362 22822
rect 4418 22820 4442 22822
rect 4202 22800 4498 22820
rect 4202 21788 4498 21808
rect 4258 21786 4282 21788
rect 4338 21786 4362 21788
rect 4418 21786 4442 21788
rect 4280 21734 4282 21786
rect 4344 21734 4356 21786
rect 4418 21734 4420 21786
rect 4258 21732 4282 21734
rect 4338 21732 4362 21734
rect 4418 21732 4442 21734
rect 4202 21712 4498 21732
rect 4202 20700 4498 20720
rect 4258 20698 4282 20700
rect 4338 20698 4362 20700
rect 4418 20698 4442 20700
rect 4280 20646 4282 20698
rect 4344 20646 4356 20698
rect 4418 20646 4420 20698
rect 4258 20644 4282 20646
rect 4338 20644 4362 20646
rect 4418 20644 4442 20646
rect 4202 20624 4498 20644
rect 4202 19612 4498 19632
rect 4258 19610 4282 19612
rect 4338 19610 4362 19612
rect 4418 19610 4442 19612
rect 4280 19558 4282 19610
rect 4344 19558 4356 19610
rect 4418 19558 4420 19610
rect 4258 19556 4282 19558
rect 4338 19556 4362 19558
rect 4418 19556 4442 19558
rect 4202 19536 4498 19556
rect 4202 18524 4498 18544
rect 4258 18522 4282 18524
rect 4338 18522 4362 18524
rect 4418 18522 4442 18524
rect 4280 18470 4282 18522
rect 4344 18470 4356 18522
rect 4418 18470 4420 18522
rect 4258 18468 4282 18470
rect 4338 18468 4362 18470
rect 4418 18468 4442 18470
rect 4202 18448 4498 18468
rect 4202 17436 4498 17456
rect 4258 17434 4282 17436
rect 4338 17434 4362 17436
rect 4418 17434 4442 17436
rect 4280 17382 4282 17434
rect 4344 17382 4356 17434
rect 4418 17382 4420 17434
rect 4258 17380 4282 17382
rect 4338 17380 4362 17382
rect 4418 17380 4442 17382
rect 4202 17360 4498 17380
rect 4202 16348 4498 16368
rect 4258 16346 4282 16348
rect 4338 16346 4362 16348
rect 4418 16346 4442 16348
rect 4280 16294 4282 16346
rect 4344 16294 4356 16346
rect 4418 16294 4420 16346
rect 4258 16292 4282 16294
rect 4338 16292 4362 16294
rect 4418 16292 4442 16294
rect 4202 16272 4498 16292
rect 4202 15260 4498 15280
rect 4258 15258 4282 15260
rect 4338 15258 4362 15260
rect 4418 15258 4442 15260
rect 4280 15206 4282 15258
rect 4344 15206 4356 15258
rect 4418 15206 4420 15258
rect 4258 15204 4282 15206
rect 4338 15204 4362 15206
rect 4418 15204 4442 15206
rect 4202 15184 4498 15204
rect 4202 14172 4498 14192
rect 4258 14170 4282 14172
rect 4338 14170 4362 14172
rect 4418 14170 4442 14172
rect 4280 14118 4282 14170
rect 4344 14118 4356 14170
rect 4418 14118 4420 14170
rect 4258 14116 4282 14118
rect 4338 14116 4362 14118
rect 4418 14116 4442 14118
rect 4202 14096 4498 14116
rect 4202 13084 4498 13104
rect 4258 13082 4282 13084
rect 4338 13082 4362 13084
rect 4418 13082 4442 13084
rect 4280 13030 4282 13082
rect 4344 13030 4356 13082
rect 4418 13030 4420 13082
rect 4258 13028 4282 13030
rect 4338 13028 4362 13030
rect 4418 13028 4442 13030
rect 4202 13008 4498 13028
rect 4202 11996 4498 12016
rect 4258 11994 4282 11996
rect 4338 11994 4362 11996
rect 4418 11994 4442 11996
rect 4280 11942 4282 11994
rect 4344 11942 4356 11994
rect 4418 11942 4420 11994
rect 4258 11940 4282 11942
rect 4338 11940 4362 11942
rect 4418 11940 4442 11942
rect 4202 11920 4498 11940
rect 4202 10908 4498 10928
rect 4258 10906 4282 10908
rect 4338 10906 4362 10908
rect 4418 10906 4442 10908
rect 4280 10854 4282 10906
rect 4344 10854 4356 10906
rect 4418 10854 4420 10906
rect 4258 10852 4282 10854
rect 4338 10852 4362 10854
rect 4418 10852 4442 10854
rect 4202 10832 4498 10852
rect 4202 9820 4498 9840
rect 4258 9818 4282 9820
rect 4338 9818 4362 9820
rect 4418 9818 4442 9820
rect 4280 9766 4282 9818
rect 4344 9766 4356 9818
rect 4418 9766 4420 9818
rect 4258 9764 4282 9766
rect 4338 9764 4362 9766
rect 4418 9764 4442 9766
rect 4202 9744 4498 9764
rect 4202 8732 4498 8752
rect 4258 8730 4282 8732
rect 4338 8730 4362 8732
rect 4418 8730 4442 8732
rect 4280 8678 4282 8730
rect 4344 8678 4356 8730
rect 4418 8678 4420 8730
rect 4258 8676 4282 8678
rect 4338 8676 4362 8678
rect 4418 8676 4442 8678
rect 4202 8656 4498 8676
rect 4202 7644 4498 7664
rect 4258 7642 4282 7644
rect 4338 7642 4362 7644
rect 4418 7642 4442 7644
rect 4280 7590 4282 7642
rect 4344 7590 4356 7642
rect 4418 7590 4420 7642
rect 4258 7588 4282 7590
rect 4338 7588 4362 7590
rect 4418 7588 4442 7590
rect 4202 7568 4498 7588
rect 4202 6556 4498 6576
rect 4258 6554 4282 6556
rect 4338 6554 4362 6556
rect 4418 6554 4442 6556
rect 4280 6502 4282 6554
rect 4344 6502 4356 6554
rect 4418 6502 4420 6554
rect 4258 6500 4282 6502
rect 4338 6500 4362 6502
rect 4418 6500 4442 6502
rect 4202 6480 4498 6500
rect 4602 5636 4654 5642
rect 4602 5578 4654 5584
rect 4202 5468 4498 5488
rect 4258 5466 4282 5468
rect 4338 5466 4362 5468
rect 4418 5466 4442 5468
rect 4280 5414 4282 5466
rect 4344 5414 4356 5466
rect 4418 5414 4420 5466
rect 4258 5412 4282 5414
rect 4338 5412 4362 5414
rect 4418 5412 4442 5414
rect 4202 5392 4498 5412
rect 4202 4380 4498 4400
rect 4258 4378 4282 4380
rect 4338 4378 4362 4380
rect 4418 4378 4442 4380
rect 4280 4326 4282 4378
rect 4344 4326 4356 4378
rect 4418 4326 4420 4378
rect 4258 4324 4282 4326
rect 4338 4324 4362 4326
rect 4418 4324 4442 4326
rect 4202 4304 4498 4324
rect 4050 4072 4102 4078
rect 4050 4014 4102 4020
rect 4202 3292 4498 3312
rect 4258 3290 4282 3292
rect 4338 3290 4362 3292
rect 4418 3290 4442 3292
rect 4280 3238 4282 3290
rect 4344 3238 4356 3290
rect 4418 3238 4420 3290
rect 4258 3236 4282 3238
rect 4338 3236 4362 3238
rect 4418 3236 4442 3238
rect 4202 3216 4498 3236
rect 4202 2204 4498 2224
rect 4258 2202 4282 2204
rect 4338 2202 4362 2204
rect 4418 2202 4442 2204
rect 4280 2150 4282 2202
rect 4344 2150 4356 2202
rect 4418 2150 4420 2202
rect 4258 2148 4282 2150
rect 4338 2148 4362 2150
rect 4418 2148 4442 2150
rect 4202 2128 4498 2148
rect 4614 1986 4642 5578
rect 4694 4140 4746 4146
rect 4694 4082 4746 4088
rect 4338 1958 4642 1986
rect 4338 800 4366 1958
rect 4706 800 4734 4082
rect 4982 4010 5010 40054
rect 5074 4078 5102 52362
rect 5442 46374 5470 59200
rect 5902 55282 5930 59200
rect 6166 59152 6218 59158
rect 6166 59094 6218 59100
rect 5890 55276 5942 55282
rect 5890 55218 5942 55224
rect 5430 46368 5482 46374
rect 5430 46310 5482 46316
rect 5154 44260 5206 44266
rect 5154 44202 5206 44208
rect 5166 4146 5194 44202
rect 5246 39296 5298 39302
rect 5246 39238 5298 39244
rect 5154 4140 5206 4146
rect 5154 4082 5206 4088
rect 5062 4072 5114 4078
rect 5062 4014 5114 4020
rect 4970 4004 5022 4010
rect 4970 3946 5022 3952
rect 5258 2666 5286 39238
rect 5614 19848 5666 19854
rect 5614 19790 5666 19796
rect 5626 19514 5654 19790
rect 5614 19508 5666 19514
rect 5614 19450 5666 19456
rect 5796 12064 5852 12073
rect 5796 11999 5852 12008
rect 5338 6656 5390 6662
rect 5338 6598 5390 6604
rect 5350 3534 5378 6598
rect 5430 4072 5482 4078
rect 5430 4014 5482 4020
rect 5338 3528 5390 3534
rect 5338 3470 5390 3476
rect 5074 2638 5286 2666
rect 5074 800 5102 2638
rect 5442 800 5470 4014
rect 5810 800 5838 11999
rect 6178 9722 6206 59094
rect 6454 55350 6482 59200
rect 6258 55344 6310 55350
rect 6258 55286 6310 55292
rect 6442 55344 6494 55350
rect 6442 55286 6494 55292
rect 6166 9716 6218 9722
rect 6166 9658 6218 9664
rect 6074 9648 6126 9654
rect 6074 9590 6126 9596
rect 6086 3194 6114 9590
rect 6166 4140 6218 4146
rect 6166 4082 6218 4088
rect 6074 3188 6126 3194
rect 6074 3130 6126 3136
rect 6178 800 6206 4082
rect 6270 3942 6298 55286
rect 7006 55282 7034 59200
rect 7270 55752 7322 55758
rect 7270 55694 7322 55700
rect 6810 55276 6862 55282
rect 6810 55218 6862 55224
rect 6994 55276 7046 55282
rect 6994 55218 7046 55224
rect 6822 37262 6850 55218
rect 6810 37256 6862 37262
rect 6810 37198 6862 37204
rect 6350 36032 6402 36038
rect 6350 35974 6402 35980
rect 6258 3936 6310 3942
rect 6258 3878 6310 3884
rect 6362 3602 6390 35974
rect 6810 26444 6862 26450
rect 6810 26386 6862 26392
rect 6718 24064 6770 24070
rect 6718 24006 6770 24012
rect 6442 12232 6494 12238
rect 6730 12186 6758 24006
rect 6822 12238 6850 26386
rect 7282 19310 7310 55694
rect 7558 52442 7586 59200
rect 8098 55888 8150 55894
rect 8098 55830 8150 55836
rect 8006 55276 8058 55282
rect 8006 55218 8058 55224
rect 7466 52414 7586 52442
rect 7466 45626 7494 52414
rect 7638 52352 7690 52358
rect 7638 52294 7690 52300
rect 7454 45620 7506 45626
rect 7454 45562 7506 45568
rect 7650 44146 7678 52294
rect 7730 45620 7782 45626
rect 7730 45562 7782 45568
rect 7914 45620 7966 45626
rect 7914 45562 7966 45568
rect 7558 44118 7678 44146
rect 7558 39370 7586 44118
rect 7362 39364 7414 39370
rect 7362 39306 7414 39312
rect 7546 39364 7598 39370
rect 7546 39306 7598 39312
rect 7374 34542 7402 39306
rect 7362 34536 7414 34542
rect 7362 34478 7414 34484
rect 7638 34536 7690 34542
rect 7638 34478 7690 34484
rect 7650 24954 7678 34478
rect 7742 29714 7770 45562
rect 7730 29708 7782 29714
rect 7730 29650 7782 29656
rect 7822 26784 7874 26790
rect 7822 26726 7874 26732
rect 7638 24948 7690 24954
rect 7638 24890 7690 24896
rect 7546 24880 7598 24886
rect 7546 24822 7598 24828
rect 7270 19304 7322 19310
rect 7270 19246 7322 19252
rect 7270 18692 7322 18698
rect 7270 18634 7322 18640
rect 7282 18426 7310 18634
rect 7270 18420 7322 18426
rect 7270 18362 7322 18368
rect 6994 14408 7046 14414
rect 6994 14350 7046 14356
rect 7006 14074 7034 14350
rect 6994 14068 7046 14074
rect 6994 14010 7046 14016
rect 6442 12174 6494 12180
rect 6454 11762 6482 12174
rect 6638 12158 6758 12186
rect 6810 12232 6862 12238
rect 6810 12174 6862 12180
rect 6442 11756 6494 11762
rect 6442 11698 6494 11704
rect 6638 7562 6666 12158
rect 6810 12096 6862 12102
rect 6808 12064 6810 12073
rect 6862 12064 6864 12073
rect 6808 11999 6864 12008
rect 6810 11756 6862 11762
rect 6810 11698 6862 11704
rect 6638 7534 6758 7562
rect 6730 4146 6758 7534
rect 6718 4140 6770 4146
rect 6718 4082 6770 4088
rect 6822 4026 6850 11698
rect 7558 9518 7586 24822
rect 7638 24200 7690 24206
rect 7638 24142 7690 24148
rect 7650 23866 7678 24142
rect 7638 23860 7690 23866
rect 7638 23802 7690 23808
rect 7834 17218 7862 26726
rect 7742 17190 7862 17218
rect 7638 14340 7690 14346
rect 7638 14282 7690 14288
rect 7546 9512 7598 9518
rect 7546 9454 7598 9460
rect 7454 4480 7506 4486
rect 7454 4422 7506 4428
rect 7466 4282 7494 4422
rect 7454 4276 7506 4282
rect 7454 4218 7506 4224
rect 7650 4146 7678 14282
rect 7742 9654 7770 17190
rect 7822 17128 7874 17134
rect 7822 17070 7874 17076
rect 7834 12306 7862 17070
rect 7822 12300 7874 12306
rect 7822 12242 7874 12248
rect 7730 9648 7782 9654
rect 7730 9590 7782 9596
rect 7730 9512 7782 9518
rect 7730 9454 7782 9460
rect 7638 4140 7690 4146
rect 7638 4082 7690 4088
rect 7742 4049 7770 9454
rect 6546 3998 6850 4026
rect 7728 4040 7784 4049
rect 6902 4004 6954 4010
rect 6350 3596 6402 3602
rect 6350 3538 6402 3544
rect 6546 800 6574 3998
rect 7728 3975 7784 3984
rect 6902 3946 6954 3952
rect 6914 800 6942 3946
rect 7270 3664 7322 3670
rect 7270 3606 7322 3612
rect 7282 800 7310 3606
rect 7926 2972 7954 45562
rect 8018 17338 8046 55218
rect 8006 17332 8058 17338
rect 8006 17274 8058 17280
rect 8006 13864 8058 13870
rect 8004 13832 8006 13841
rect 8058 13832 8060 13841
rect 8004 13767 8060 13776
rect 8110 13274 8138 55830
rect 8570 55826 8598 59200
rect 9122 59106 9150 59200
rect 8754 59078 9150 59106
rect 8558 55820 8610 55826
rect 8558 55762 8610 55768
rect 8190 55344 8242 55350
rect 8190 55286 8242 55292
rect 8202 26790 8230 55286
rect 8282 55276 8334 55282
rect 8282 55218 8334 55224
rect 8190 26784 8242 26790
rect 8190 26726 8242 26732
rect 8190 25696 8242 25702
rect 8190 25638 8242 25644
rect 8202 25498 8230 25638
rect 8190 25492 8242 25498
rect 8190 25434 8242 25440
rect 8294 20482 8322 55218
rect 8754 48346 8782 59078
rect 9582 55282 9610 59200
rect 10134 59106 10162 59200
rect 9950 59078 10162 59106
rect 10686 59106 10714 59200
rect 11238 59106 11266 59200
rect 10686 59078 10990 59106
rect 11238 59078 11358 59106
rect 9846 55956 9898 55962
rect 9846 55898 9898 55904
rect 9570 55276 9622 55282
rect 9570 55218 9622 55224
rect 8650 48340 8702 48346
rect 8650 48282 8702 48288
rect 8742 48340 8794 48346
rect 8742 48282 8794 48288
rect 8662 37330 8690 48282
rect 9202 45824 9254 45830
rect 9202 45766 9254 45772
rect 8650 37324 8702 37330
rect 8650 37266 8702 37272
rect 8742 37324 8794 37330
rect 8742 37266 8794 37272
rect 8754 32434 8782 37266
rect 9214 32774 9242 45766
rect 9570 45416 9622 45422
rect 9570 45358 9622 45364
rect 9202 32768 9254 32774
rect 9202 32710 9254 32716
rect 9478 32768 9530 32774
rect 9478 32710 9530 32716
rect 8742 32428 8794 32434
rect 8742 32370 8794 32376
rect 9202 32428 9254 32434
rect 9202 32370 9254 32376
rect 8742 31272 8794 31278
rect 8742 31214 8794 31220
rect 8754 30870 8782 31214
rect 8834 31136 8886 31142
rect 9018 31136 9070 31142
rect 8886 31084 9018 31090
rect 8834 31078 9070 31084
rect 8846 31062 9058 31078
rect 8742 30864 8794 30870
rect 8742 30806 8794 30812
rect 8466 30184 8518 30190
rect 8466 30126 8518 30132
rect 8478 29646 8506 30126
rect 8834 30048 8886 30054
rect 9018 30048 9070 30054
rect 8886 29996 9018 30002
rect 8834 29990 9070 29996
rect 8846 29974 9058 29990
rect 8466 29640 8518 29646
rect 8466 29582 8518 29588
rect 8834 29572 8886 29578
rect 8834 29514 8886 29520
rect 8846 29170 8874 29514
rect 8834 29164 8886 29170
rect 8834 29106 8886 29112
rect 8570 28082 8966 28098
rect 8558 28076 8978 28082
rect 8610 28070 8926 28076
rect 8558 28018 8610 28024
rect 8926 28018 8978 28024
rect 8834 28008 8886 28014
rect 8570 27956 8834 27962
rect 8570 27950 8886 27956
rect 8570 27934 8874 27950
rect 8570 27878 8598 27934
rect 8558 27872 8610 27878
rect 9214 27826 9242 32370
rect 8558 27814 8610 27820
rect 9168 27798 9242 27826
rect 9168 27554 9196 27798
rect 9490 27674 9518 32710
rect 9294 27668 9346 27674
rect 9294 27610 9346 27616
rect 9478 27668 9530 27674
rect 9478 27610 9530 27616
rect 9168 27526 9242 27554
rect 8834 27056 8886 27062
rect 8432 27028 8834 27044
rect 8420 27022 8834 27028
rect 8472 27016 8834 27022
rect 8834 26998 8886 27004
rect 8420 26964 8472 26970
rect 8558 26920 8610 26926
rect 8834 26920 8886 26926
rect 8610 26868 8834 26874
rect 8558 26862 8886 26868
rect 8570 26846 8874 26862
rect 8696 26784 8748 26790
rect 8696 26726 8748 26732
rect 8708 26586 8736 26726
rect 8696 26580 8748 26586
rect 8696 26522 8748 26528
rect 8558 25832 8610 25838
rect 8610 25780 8874 25786
rect 8558 25774 8874 25780
rect 8570 25758 8874 25774
rect 8846 25702 8874 25758
rect 8696 25696 8748 25702
rect 8696 25638 8748 25644
rect 8834 25696 8886 25702
rect 8834 25638 8886 25644
rect 8708 25430 8736 25638
rect 8696 25424 8748 25430
rect 8696 25366 8748 25372
rect 9018 24948 9070 24954
rect 8846 24920 9018 24936
rect 8834 24914 9018 24920
rect 8886 24908 9018 24914
rect 9018 24890 9070 24896
rect 8834 24856 8886 24862
rect 8604 24710 8656 24716
rect 8466 24676 8518 24682
rect 9018 24676 9070 24682
rect 8656 24658 9018 24664
rect 8604 24652 9018 24658
rect 8616 24636 9018 24652
rect 8466 24618 8518 24624
rect 9018 24618 9070 24624
rect 8478 24410 8506 24618
rect 8466 24404 8518 24410
rect 8466 24346 8518 24352
rect 8662 23866 8874 23882
rect 8650 23860 8886 23866
rect 8702 23854 8834 23860
rect 8650 23802 8702 23808
rect 8834 23802 8886 23808
rect 8420 23622 8472 23628
rect 8472 23594 8782 23610
rect 8472 23588 8794 23594
rect 8472 23582 8742 23588
rect 8420 23564 8472 23570
rect 8742 23530 8794 23536
rect 8466 21344 8518 21350
rect 8650 21344 8702 21350
rect 8518 21292 8650 21298
rect 8466 21286 8702 21292
rect 8478 21270 8690 21286
rect 8466 20596 8518 20602
rect 8518 20556 8598 20584
rect 8466 20538 8518 20544
rect 8294 20454 8368 20482
rect 8340 20210 8368 20454
rect 8420 20358 8472 20364
rect 8420 20300 8472 20306
rect 8294 20182 8368 20210
rect 8190 19168 8242 19174
rect 8188 19136 8190 19145
rect 8242 19136 8244 19145
rect 8188 19071 8244 19080
rect 8110 13246 8184 13274
rect 8156 12986 8184 13246
rect 8144 12980 8196 12986
rect 8144 12922 8196 12928
rect 8096 11792 8152 11801
rect 8096 11727 8098 11736
rect 8150 11727 8152 11736
rect 8098 11698 8150 11704
rect 8098 9648 8150 9654
rect 8098 9590 8150 9596
rect 8110 4146 8138 9590
rect 8190 6724 8242 6730
rect 8190 6666 8242 6672
rect 8202 6458 8230 6666
rect 8190 6452 8242 6458
rect 8190 6394 8242 6400
rect 8294 6338 8322 20182
rect 8432 20074 8460 20300
rect 8432 20058 8506 20074
rect 8432 20052 8518 20058
rect 8432 20046 8466 20052
rect 8466 19994 8518 20000
rect 8466 19508 8518 19514
rect 8466 19450 8518 19456
rect 8478 19417 8506 19450
rect 8464 19408 8520 19417
rect 8464 19343 8520 19352
rect 8420 19270 8472 19276
rect 8420 19212 8472 19218
rect 8432 18986 8460 19212
rect 8432 18970 8506 18986
rect 8432 18964 8518 18970
rect 8432 18958 8466 18964
rect 8466 18906 8518 18912
rect 8570 18902 8598 20556
rect 8926 19168 8978 19174
rect 8924 19136 8926 19145
rect 8978 19136 8980 19145
rect 8924 19071 8980 19080
rect 8558 18896 8610 18902
rect 8558 18838 8610 18844
rect 8846 18426 9058 18442
rect 8834 18420 9070 18426
rect 8886 18414 9018 18420
rect 8834 18362 8886 18368
rect 9018 18362 9070 18368
rect 9214 18034 9242 27526
rect 9168 18006 9242 18034
rect 9168 17898 9196 18006
rect 9122 17870 9196 17898
rect 8834 17808 8886 17814
rect 8834 17750 8886 17756
rect 8742 17740 8794 17746
rect 8742 17682 8794 17688
rect 8754 17134 8782 17682
rect 8846 17338 8874 17750
rect 8834 17332 8886 17338
rect 8834 17274 8886 17280
rect 8742 17128 8794 17134
rect 8742 17070 8794 17076
rect 8650 16448 8702 16454
rect 8650 16390 8702 16396
rect 8662 16132 8690 16390
rect 8742 16244 8794 16250
rect 8742 16186 8794 16192
rect 8650 16126 8702 16132
rect 8650 16068 8702 16074
rect 8754 15910 8782 16186
rect 8742 15904 8794 15910
rect 8742 15846 8794 15852
rect 8478 15162 8690 15178
rect 8466 15156 8702 15162
rect 8518 15150 8650 15156
rect 8466 15098 8518 15104
rect 8650 15098 8702 15104
rect 8650 15020 8702 15026
rect 8650 14962 8702 14968
rect 8374 14918 8426 14924
rect 8662 14906 8690 14962
rect 8426 14878 8690 14906
rect 8374 14860 8426 14866
rect 8374 9478 8426 9484
rect 8374 9420 8426 9426
rect 8386 9178 8414 9420
rect 8374 9172 8426 9178
rect 8374 9114 8426 9120
rect 8570 8498 8874 8514
rect 8570 8492 8886 8498
rect 8570 8486 8834 8492
rect 8570 8430 8598 8486
rect 8834 8434 8886 8440
rect 8558 8424 8610 8430
rect 8558 8366 8610 8372
rect 8386 7410 8690 7426
rect 8386 7404 8702 7410
rect 8386 7398 8650 7404
rect 8386 7342 8414 7398
rect 8650 7346 8702 7352
rect 8374 7336 8426 7342
rect 8374 7278 8426 7284
rect 8466 6656 8518 6662
rect 8466 6598 8518 6604
rect 8478 6458 8506 6598
rect 8466 6452 8518 6458
rect 8466 6394 8518 6400
rect 8294 6310 8368 6338
rect 8340 6066 8368 6310
rect 8340 6038 8414 6066
rect 8236 5262 8288 5268
rect 8386 5250 8414 6038
rect 8466 5908 8518 5914
rect 8466 5850 8518 5856
rect 8288 5222 8414 5250
rect 8236 5204 8288 5210
rect 8006 4140 8058 4146
rect 8006 4082 8058 4088
rect 8098 4140 8150 4146
rect 8098 4082 8150 4088
rect 7650 2944 7954 2972
rect 7650 800 7678 2944
rect 8018 800 8046 4082
rect 8374 3732 8426 3738
rect 8374 3674 8426 3680
rect 8386 800 8414 3674
rect 8478 3058 8506 5850
rect 8742 5160 8794 5166
rect 8742 5102 8794 5108
rect 8650 5024 8702 5030
rect 8754 4978 8782 5102
rect 8702 4972 8782 4978
rect 8650 4966 8782 4972
rect 8662 4950 8782 4966
rect 9122 4282 9150 17870
rect 9202 17298 9254 17304
rect 9202 17241 9254 17246
rect 9200 17232 9256 17241
rect 9200 17167 9256 17176
rect 9306 13682 9334 27610
rect 9478 20460 9530 20466
rect 9478 20402 9530 20408
rect 9214 13654 9334 13682
rect 9110 4276 9162 4282
rect 9110 4218 9162 4224
rect 8834 3120 8886 3126
rect 9214 3097 9242 13654
rect 9490 13138 9518 20402
rect 9398 13110 9518 13138
rect 9294 11008 9346 11014
rect 9294 10950 9346 10956
rect 9306 10538 9334 10950
rect 9294 10532 9346 10538
rect 9294 10474 9346 10480
rect 8834 3062 8886 3068
rect 9200 3088 9256 3097
rect 8466 3052 8518 3058
rect 8466 2994 8518 3000
rect 8846 1714 8874 3062
rect 9200 3023 9256 3032
rect 9398 2938 9426 13110
rect 9582 7562 9610 45358
rect 9858 10606 9886 55898
rect 9950 42226 9978 59078
rect 10858 56364 10910 56370
rect 10858 56306 10910 56312
rect 10582 56296 10634 56302
rect 10582 56238 10634 56244
rect 10490 55684 10542 55690
rect 10490 55626 10542 55632
rect 10306 46980 10358 46986
rect 10306 46922 10358 46928
rect 9938 42220 9990 42226
rect 9938 42162 9990 42168
rect 10318 22794 10346 46922
rect 10042 22766 10346 22794
rect 9662 10600 9714 10606
rect 9662 10542 9714 10548
rect 9846 10600 9898 10606
rect 9846 10542 9898 10548
rect 9674 10266 9702 10542
rect 9662 10260 9714 10266
rect 9662 10202 9714 10208
rect 8754 1686 8874 1714
rect 9122 2910 9426 2938
rect 9490 7534 9610 7562
rect 8754 800 8782 1686
rect 9122 800 9150 2910
rect 9490 800 9518 7534
rect 10042 6730 10070 22766
rect 10398 18964 10450 18970
rect 10398 18906 10450 18912
rect 10410 9994 10438 18906
rect 10398 9988 10450 9994
rect 10398 9930 10450 9936
rect 10502 9874 10530 55626
rect 10594 46986 10622 56238
rect 10870 51474 10898 56306
rect 10858 51468 10910 51474
rect 10858 51410 10910 51416
rect 10582 46980 10634 46986
rect 10582 46922 10634 46928
rect 10858 20392 10910 20398
rect 10858 20334 10910 20340
rect 10582 14068 10634 14074
rect 10582 14010 10634 14016
rect 10134 9846 10530 9874
rect 10030 6724 10082 6730
rect 10030 6666 10082 6672
rect 10134 6662 10162 9846
rect 10594 9738 10622 14010
rect 10766 12776 10818 12782
rect 10766 12718 10818 12724
rect 10674 9988 10726 9994
rect 10674 9930 10726 9936
rect 10226 9710 10622 9738
rect 10122 6656 10174 6662
rect 10122 6598 10174 6604
rect 9846 4140 9898 4146
rect 9846 4082 9898 4088
rect 9570 2848 9622 2854
rect 9570 2790 9622 2796
rect 9582 2514 9610 2790
rect 9570 2508 9622 2514
rect 9570 2450 9622 2456
rect 9858 800 9886 4082
rect 10226 800 10254 9710
rect 10582 6248 10634 6254
rect 10582 6190 10634 6196
rect 10594 800 10622 6190
rect 10686 3942 10714 9930
rect 10778 4146 10806 12718
rect 10870 9654 10898 20334
rect 10962 19786 10990 59078
rect 11134 37120 11186 37126
rect 11134 37062 11186 37068
rect 11042 31272 11094 31278
rect 11042 31214 11094 31220
rect 11054 30938 11082 31214
rect 11042 30932 11094 30938
rect 11042 30874 11094 30880
rect 10950 19780 11002 19786
rect 10950 19722 11002 19728
rect 10858 9648 10910 9654
rect 10858 9590 10910 9596
rect 10858 9512 10910 9518
rect 10858 9454 10910 9460
rect 11042 9512 11094 9518
rect 11042 9454 11094 9460
rect 10766 4140 10818 4146
rect 10766 4082 10818 4088
rect 10674 3936 10726 3942
rect 10674 3878 10726 3884
rect 10870 3194 10898 9454
rect 10950 8356 11002 8362
rect 10950 8298 11002 8304
rect 10858 3188 10910 3194
rect 10858 3130 10910 3136
rect 10962 800 10990 8298
rect 11054 3670 11082 9454
rect 11042 3664 11094 3670
rect 11146 3641 11174 37062
rect 11226 31272 11278 31278
rect 11226 31214 11278 31220
rect 11042 3606 11094 3612
rect 11132 3632 11188 3641
rect 11132 3567 11188 3576
rect 11238 3505 11266 31214
rect 11330 5234 11358 59078
rect 11698 55282 11726 59200
rect 11686 55276 11738 55282
rect 11686 55218 11738 55224
rect 12146 55276 12198 55282
rect 12146 55218 12198 55224
rect 11778 36712 11830 36718
rect 11778 36654 11830 36660
rect 11502 18216 11554 18222
rect 11502 18158 11554 18164
rect 11514 12374 11542 18158
rect 11502 12368 11554 12374
rect 11502 12310 11554 12316
rect 11686 11892 11738 11898
rect 11686 11834 11738 11840
rect 11698 11801 11726 11834
rect 11684 11792 11740 11801
rect 11684 11727 11740 11736
rect 11318 5228 11370 5234
rect 11318 5170 11370 5176
rect 11686 4140 11738 4146
rect 11686 4082 11738 4088
rect 11318 4072 11370 4078
rect 11318 4014 11370 4020
rect 11224 3496 11280 3505
rect 11224 3431 11280 3440
rect 11330 800 11358 4014
rect 11698 800 11726 4082
rect 11790 3738 11818 36654
rect 11870 32768 11922 32774
rect 11870 32710 11922 32716
rect 11882 32570 11910 32710
rect 11870 32564 11922 32570
rect 11870 32506 11922 32512
rect 12054 29096 12106 29102
rect 12054 29038 12106 29044
rect 11870 9648 11922 9654
rect 11870 9590 11922 9596
rect 11882 3738 11910 9590
rect 12066 4078 12094 29038
rect 12158 26382 12186 55218
rect 12146 26376 12198 26382
rect 12146 26318 12198 26324
rect 12250 7818 12278 59200
rect 12802 55162 12830 59200
rect 13066 55820 13118 55826
rect 13066 55762 13118 55768
rect 12434 55134 12830 55162
rect 12330 53032 12382 53038
rect 12330 52974 12382 52980
rect 12238 7812 12290 7818
rect 12238 7754 12290 7760
rect 12342 4146 12370 52974
rect 12434 5370 12462 55134
rect 12790 24132 12842 24138
rect 12790 24074 12842 24080
rect 12802 23662 12830 24074
rect 13078 23798 13106 55762
rect 13262 55622 13290 59200
rect 13618 56500 13670 56506
rect 13618 56442 13670 56448
rect 13250 55616 13302 55622
rect 13250 55558 13302 55564
rect 13526 42152 13578 42158
rect 13526 42094 13578 42100
rect 13158 30184 13210 30190
rect 13158 30126 13210 30132
rect 13170 29850 13198 30126
rect 13158 29844 13210 29850
rect 13158 29786 13210 29792
rect 13342 27668 13394 27674
rect 13342 27610 13394 27616
rect 12882 23792 12934 23798
rect 12882 23734 12934 23740
rect 13066 23792 13118 23798
rect 13066 23734 13118 23740
rect 12790 23656 12842 23662
rect 12790 23598 12842 23604
rect 12894 23594 12922 23734
rect 12882 23588 12934 23594
rect 12882 23530 12934 23536
rect 13066 19168 13118 19174
rect 13066 19110 13118 19116
rect 12790 18080 12842 18086
rect 12790 18022 12842 18028
rect 12514 13864 12566 13870
rect 12512 13832 12514 13841
rect 12566 13832 12568 13841
rect 12512 13767 12568 13776
rect 12422 5364 12474 5370
rect 12422 5306 12474 5312
rect 12802 4826 12830 18022
rect 13078 7698 13106 19110
rect 13354 12458 13382 27610
rect 13434 21888 13486 21894
rect 13434 21830 13486 21836
rect 12894 7670 13106 7698
rect 13170 12430 13382 12458
rect 12790 4820 12842 4826
rect 12790 4762 12842 4768
rect 12330 4140 12382 4146
rect 12330 4082 12382 4088
rect 12054 4072 12106 4078
rect 12054 4014 12106 4020
rect 12790 4004 12842 4010
rect 12790 3946 12842 3952
rect 11778 3732 11830 3738
rect 11778 3674 11830 3680
rect 11870 3732 11922 3738
rect 11870 3674 11922 3680
rect 12054 2848 12106 2854
rect 12054 2790 12106 2796
rect 12066 800 12094 2790
rect 12422 2508 12474 2514
rect 12422 2450 12474 2456
rect 12434 800 12462 2450
rect 12802 800 12830 3946
rect 12894 3670 12922 7670
rect 12974 4820 13026 4826
rect 12974 4762 13026 4768
rect 12882 3664 12934 3670
rect 12882 3606 12934 3612
rect 12986 800 13014 4762
rect 13066 4140 13118 4146
rect 13066 4082 13118 4088
rect 13078 800 13106 4082
rect 13170 2514 13198 12430
rect 13250 12368 13302 12374
rect 13250 12310 13302 12316
rect 13262 4026 13290 12310
rect 13446 4298 13474 21830
rect 13354 4270 13474 4298
rect 13354 4146 13382 4270
rect 13342 4140 13394 4146
rect 13342 4082 13394 4088
rect 13434 4140 13486 4146
rect 13434 4082 13486 4088
rect 13262 3998 13382 4026
rect 13158 2508 13210 2514
rect 13158 2450 13210 2456
rect 13354 800 13382 3998
rect 13446 800 13474 4082
rect 13538 4010 13566 42094
rect 13630 26042 13658 56442
rect 13814 55282 13842 59200
rect 14446 56432 14498 56438
rect 14446 56374 14498 56380
rect 13802 55276 13854 55282
rect 13802 55218 13854 55224
rect 13802 51060 13854 51066
rect 13802 51002 13854 51008
rect 13710 48680 13762 48686
rect 13710 48622 13762 48628
rect 13618 26036 13670 26042
rect 13618 25978 13670 25984
rect 13618 18284 13670 18290
rect 13618 18226 13670 18232
rect 13526 4004 13578 4010
rect 13526 3946 13578 3952
rect 13630 2802 13658 18226
rect 13722 4146 13750 48622
rect 13814 15094 13842 51002
rect 13894 28212 13946 28218
rect 13894 28154 13946 28160
rect 13906 27674 13934 28154
rect 13894 27668 13946 27674
rect 13894 27610 13946 27616
rect 14170 18420 14222 18426
rect 14170 18362 14222 18368
rect 13802 15088 13854 15094
rect 13802 15030 13854 15036
rect 13710 4140 13762 4146
rect 13710 4082 13762 4088
rect 13802 4072 13854 4078
rect 13802 4014 13854 4020
rect 13538 2774 13658 2802
rect 13538 2666 13566 2774
rect 13538 2638 13750 2666
rect 13722 800 13750 2638
rect 13814 800 13842 4014
rect 14182 800 14210 18362
rect 14458 6118 14486 56374
rect 14918 51066 14946 59200
rect 14998 55344 15050 55350
rect 14998 55286 15050 55292
rect 14906 51060 14958 51066
rect 14906 51002 14958 51008
rect 15010 43450 15038 55286
rect 15090 55276 15142 55282
rect 15090 55218 15142 55224
rect 14998 43444 15050 43450
rect 14998 43386 15050 43392
rect 14630 40112 14682 40118
rect 14630 40054 14682 40060
rect 14538 20256 14590 20262
rect 14538 20198 14590 20204
rect 14446 6112 14498 6118
rect 14446 6054 14498 6060
rect 14550 4146 14578 20198
rect 14538 4140 14590 4146
rect 14538 4082 14590 4088
rect 14446 3936 14498 3942
rect 14446 3878 14498 3884
rect 14352 3768 14408 3777
rect 14352 3703 14408 3712
rect 14366 3602 14394 3703
rect 14354 3596 14406 3602
rect 14354 3538 14406 3544
rect 14458 800 14486 3878
rect 14642 3398 14670 40054
rect 14998 30184 15050 30190
rect 14998 30126 15050 30132
rect 14906 5568 14958 5574
rect 14906 5510 14958 5516
rect 14814 3664 14866 3670
rect 14814 3606 14866 3612
rect 14630 3392 14682 3398
rect 14630 3334 14682 3340
rect 14538 2304 14590 2310
rect 14538 2246 14590 2252
rect 14550 800 14578 2246
rect 14826 800 14854 3606
rect 14918 800 14946 5510
rect 15010 4078 15038 30126
rect 15102 16046 15130 55218
rect 15378 52714 15406 59200
rect 15826 56704 15878 56710
rect 15826 56646 15878 56652
rect 15838 56114 15866 56646
rect 15930 56302 15958 59200
rect 15918 56296 15970 56302
rect 15918 56238 15970 56244
rect 16482 56234 16510 59200
rect 16470 56228 16522 56234
rect 16470 56170 16522 56176
rect 15838 56086 15958 56114
rect 15286 52686 15406 52714
rect 15090 16040 15142 16046
rect 15090 15982 15142 15988
rect 15182 15904 15234 15910
rect 15180 15872 15182 15881
rect 15234 15872 15236 15881
rect 15180 15807 15236 15816
rect 15182 11892 15234 11898
rect 15182 11834 15234 11840
rect 15194 11801 15222 11834
rect 15180 11792 15236 11801
rect 15180 11727 15236 11736
rect 15286 5166 15314 52686
rect 15642 29504 15694 29510
rect 15642 29446 15694 29452
rect 15654 22794 15682 29446
rect 15654 22766 15774 22794
rect 15548 19408 15604 19417
rect 15548 19343 15604 19352
rect 15562 13138 15590 19343
rect 15378 13110 15590 13138
rect 15274 5160 15326 5166
rect 15274 5102 15326 5108
rect 15378 4842 15406 13110
rect 15642 7880 15694 7886
rect 15642 7822 15694 7828
rect 15286 4814 15406 4842
rect 14998 4072 15050 4078
rect 14998 4014 15050 4020
rect 15286 800 15314 4814
rect 15458 4140 15510 4146
rect 15458 4082 15510 4088
rect 15470 800 15498 4082
rect 15654 800 15682 7822
rect 15746 3942 15774 22766
rect 15930 7750 15958 56086
rect 17034 55350 17062 59200
rect 17494 55690 17522 59200
rect 18046 55758 18074 59200
rect 18492 55856 18548 55865
rect 18492 55791 18548 55800
rect 18034 55752 18086 55758
rect 18034 55694 18086 55700
rect 17482 55684 17534 55690
rect 17482 55626 17534 55632
rect 17574 55412 17626 55418
rect 17574 55354 17626 55360
rect 17022 55344 17074 55350
rect 17022 55286 17074 55292
rect 16470 49768 16522 49774
rect 16470 49710 16522 49716
rect 16378 44736 16430 44742
rect 16378 44678 16430 44684
rect 16194 20324 16246 20330
rect 16194 20266 16246 20272
rect 15918 7744 15970 7750
rect 15918 7686 15970 7692
rect 15826 7540 15878 7546
rect 15826 7482 15878 7488
rect 15734 3936 15786 3942
rect 15734 3878 15786 3884
rect 15838 800 15866 7482
rect 16010 4140 16062 4146
rect 16010 4082 16062 4088
rect 16022 800 16050 4082
rect 16206 800 16234 20266
rect 16286 20052 16338 20058
rect 16286 19994 16338 20000
rect 16298 7546 16326 19994
rect 16390 7886 16418 44678
rect 16378 7880 16430 7886
rect 16378 7822 16430 7828
rect 16378 7744 16430 7750
rect 16378 7686 16430 7692
rect 16286 7540 16338 7546
rect 16286 7482 16338 7488
rect 16286 7336 16338 7342
rect 16286 7278 16338 7284
rect 16298 3058 16326 7278
rect 16286 3052 16338 3058
rect 16286 2994 16338 3000
rect 16390 800 16418 7686
rect 16482 4146 16510 49710
rect 17586 46986 17614 55354
rect 18126 54528 18178 54534
rect 18126 54470 18178 54476
rect 17206 46980 17258 46986
rect 17206 46922 17258 46928
rect 17574 46980 17626 46986
rect 17574 46922 17626 46928
rect 16562 27056 16614 27062
rect 16562 26998 16614 27004
rect 16574 26858 16602 26998
rect 16562 26852 16614 26858
rect 16562 26794 16614 26800
rect 17218 22794 17246 46922
rect 17850 45348 17902 45354
rect 17850 45290 17902 45296
rect 17218 22766 17338 22794
rect 17022 21548 17074 21554
rect 17022 21490 17074 21496
rect 16930 21480 16982 21486
rect 16930 21422 16982 21428
rect 16838 21344 16890 21350
rect 16838 21286 16890 21292
rect 16746 18896 16798 18902
rect 16746 18838 16798 18844
rect 16470 4140 16522 4146
rect 16470 4082 16522 4088
rect 16758 800 16786 18838
rect 16850 4010 16878 21286
rect 16838 4004 16890 4010
rect 16838 3946 16890 3952
rect 16942 800 16970 21422
rect 17034 4826 17062 21490
rect 17114 13184 17166 13190
rect 17114 13126 17166 13132
rect 17126 12986 17154 13126
rect 17114 12980 17166 12986
rect 17114 12922 17166 12928
rect 17310 6458 17338 22766
rect 17482 9716 17534 9722
rect 17482 9658 17534 9664
rect 17298 6452 17350 6458
rect 17298 6394 17350 6400
rect 17022 4820 17074 4826
rect 17022 4762 17074 4768
rect 17390 4820 17442 4826
rect 17390 4762 17442 4768
rect 17114 4140 17166 4146
rect 17114 4082 17166 4088
rect 17126 800 17154 4082
rect 17298 3596 17350 3602
rect 17298 3538 17350 3544
rect 17310 3194 17338 3538
rect 17298 3188 17350 3194
rect 17298 3130 17350 3136
rect 17402 898 17430 4762
rect 17310 870 17430 898
rect 17310 800 17338 870
rect 17494 800 17522 9658
rect 17862 4146 17890 45290
rect 18034 22500 18086 22506
rect 18034 22442 18086 22448
rect 17942 18692 17994 18698
rect 17942 18634 17994 18640
rect 17850 4140 17902 4146
rect 17850 4082 17902 4088
rect 17850 4004 17902 4010
rect 17850 3946 17902 3952
rect 17862 800 17890 3946
rect 17954 1426 17982 18634
rect 17942 1420 17994 1426
rect 17942 1362 17994 1368
rect 18046 800 18074 22442
rect 18138 3369 18166 54470
rect 18506 53394 18534 55791
rect 18598 55282 18626 59200
rect 18678 55684 18730 55690
rect 18678 55626 18730 55632
rect 18586 55276 18638 55282
rect 18586 55218 18638 55224
rect 18506 53366 18626 53394
rect 18218 50856 18270 50862
rect 18218 50798 18270 50804
rect 18124 3360 18180 3369
rect 18124 3295 18180 3304
rect 18230 3233 18258 50798
rect 18402 22772 18454 22778
rect 18402 22714 18454 22720
rect 18310 22568 18362 22574
rect 18310 22510 18362 22516
rect 18322 7546 18350 22510
rect 18414 14550 18442 22714
rect 18494 22432 18546 22438
rect 18494 22374 18546 22380
rect 18402 14544 18454 14550
rect 18402 14486 18454 14492
rect 18310 7540 18362 7546
rect 18310 7482 18362 7488
rect 18506 4842 18534 22374
rect 18414 4814 18534 4842
rect 18216 3224 18272 3233
rect 18216 3159 18272 3168
rect 18218 1420 18270 1426
rect 18218 1362 18270 1368
rect 18230 800 18258 1362
rect 18414 800 18442 4814
rect 18598 3194 18626 53366
rect 18690 15094 18718 55626
rect 19058 49178 19086 59200
rect 19610 57338 19638 59200
rect 19610 57310 19914 57338
rect 19562 57148 19858 57168
rect 19618 57146 19642 57148
rect 19698 57146 19722 57148
rect 19778 57146 19802 57148
rect 19640 57094 19642 57146
rect 19704 57094 19716 57146
rect 19778 57094 19780 57146
rect 19618 57092 19642 57094
rect 19698 57092 19722 57094
rect 19778 57092 19802 57094
rect 19562 57072 19858 57092
rect 19562 56060 19858 56080
rect 19618 56058 19642 56060
rect 19698 56058 19722 56060
rect 19778 56058 19802 56060
rect 19640 56006 19642 56058
rect 19704 56006 19716 56058
rect 19778 56006 19780 56058
rect 19618 56004 19642 56006
rect 19698 56004 19722 56006
rect 19778 56004 19802 56006
rect 19562 55984 19858 56004
rect 19414 55752 19466 55758
rect 19414 55694 19466 55700
rect 19138 55276 19190 55282
rect 19138 55218 19190 55224
rect 18782 49150 19086 49178
rect 18782 37346 18810 49150
rect 18862 49088 18914 49094
rect 18862 49030 18914 49036
rect 18874 48346 18902 49030
rect 18862 48340 18914 48346
rect 18862 48282 18914 48288
rect 18954 48340 19006 48346
rect 18954 48282 19006 48288
rect 18966 38570 18994 48282
rect 19150 39098 19178 55218
rect 19320 54632 19376 54641
rect 19320 54567 19322 54576
rect 19374 54567 19376 54576
rect 19322 54538 19374 54544
rect 19138 39092 19190 39098
rect 19138 39034 19190 39040
rect 18966 38542 19178 38570
rect 18782 37318 18902 37346
rect 18874 29073 18902 37318
rect 18860 29064 18916 29073
rect 19150 29034 19178 38542
rect 19426 36922 19454 55694
rect 19886 55282 19914 57310
rect 19966 56296 20018 56302
rect 19966 56238 20018 56244
rect 19874 55276 19926 55282
rect 19874 55218 19926 55224
rect 19562 54972 19858 54992
rect 19618 54970 19642 54972
rect 19698 54970 19722 54972
rect 19778 54970 19802 54972
rect 19640 54918 19642 54970
rect 19704 54918 19716 54970
rect 19778 54918 19780 54970
rect 19618 54916 19642 54918
rect 19698 54916 19722 54918
rect 19778 54916 19802 54918
rect 19562 54896 19858 54916
rect 19562 53884 19858 53904
rect 19618 53882 19642 53884
rect 19698 53882 19722 53884
rect 19778 53882 19802 53884
rect 19640 53830 19642 53882
rect 19704 53830 19716 53882
rect 19778 53830 19780 53882
rect 19618 53828 19642 53830
rect 19698 53828 19722 53830
rect 19778 53828 19802 53830
rect 19562 53808 19858 53828
rect 19978 53666 20006 56238
rect 20162 55978 20190 59200
rect 20162 55950 20558 55978
rect 20150 55820 20202 55826
rect 20150 55762 20202 55768
rect 20058 55344 20110 55350
rect 20058 55286 20110 55292
rect 19886 53638 20006 53666
rect 19562 52796 19858 52816
rect 19618 52794 19642 52796
rect 19698 52794 19722 52796
rect 19778 52794 19802 52796
rect 19640 52742 19642 52794
rect 19704 52742 19716 52794
rect 19778 52742 19780 52794
rect 19618 52740 19642 52742
rect 19698 52740 19722 52742
rect 19778 52740 19802 52742
rect 19562 52720 19858 52740
rect 19562 51708 19858 51728
rect 19618 51706 19642 51708
rect 19698 51706 19722 51708
rect 19778 51706 19802 51708
rect 19640 51654 19642 51706
rect 19704 51654 19716 51706
rect 19778 51654 19780 51706
rect 19618 51652 19642 51654
rect 19698 51652 19722 51654
rect 19778 51652 19802 51654
rect 19562 51632 19858 51652
rect 19562 50620 19858 50640
rect 19618 50618 19642 50620
rect 19698 50618 19722 50620
rect 19778 50618 19802 50620
rect 19640 50566 19642 50618
rect 19704 50566 19716 50618
rect 19778 50566 19780 50618
rect 19618 50564 19642 50566
rect 19698 50564 19722 50566
rect 19778 50564 19802 50566
rect 19562 50544 19858 50564
rect 19562 49532 19858 49552
rect 19618 49530 19642 49532
rect 19698 49530 19722 49532
rect 19778 49530 19802 49532
rect 19640 49478 19642 49530
rect 19704 49478 19716 49530
rect 19778 49478 19780 49530
rect 19618 49476 19642 49478
rect 19698 49476 19722 49478
rect 19778 49476 19802 49478
rect 19562 49456 19858 49476
rect 19562 48444 19858 48464
rect 19618 48442 19642 48444
rect 19698 48442 19722 48444
rect 19778 48442 19802 48444
rect 19640 48390 19642 48442
rect 19704 48390 19716 48442
rect 19778 48390 19780 48442
rect 19618 48388 19642 48390
rect 19698 48388 19722 48390
rect 19778 48388 19802 48390
rect 19562 48368 19858 48388
rect 19562 47356 19858 47376
rect 19618 47354 19642 47356
rect 19698 47354 19722 47356
rect 19778 47354 19802 47356
rect 19640 47302 19642 47354
rect 19704 47302 19716 47354
rect 19778 47302 19780 47354
rect 19618 47300 19642 47302
rect 19698 47300 19722 47302
rect 19778 47300 19802 47302
rect 19562 47280 19858 47300
rect 19562 46268 19858 46288
rect 19618 46266 19642 46268
rect 19698 46266 19722 46268
rect 19778 46266 19802 46268
rect 19640 46214 19642 46266
rect 19704 46214 19716 46266
rect 19778 46214 19780 46266
rect 19618 46212 19642 46214
rect 19698 46212 19722 46214
rect 19778 46212 19802 46214
rect 19562 46192 19858 46212
rect 19562 45180 19858 45200
rect 19618 45178 19642 45180
rect 19698 45178 19722 45180
rect 19778 45178 19802 45180
rect 19640 45126 19642 45178
rect 19704 45126 19716 45178
rect 19778 45126 19780 45178
rect 19618 45124 19642 45126
rect 19698 45124 19722 45126
rect 19778 45124 19802 45126
rect 19562 45104 19858 45124
rect 19562 44092 19858 44112
rect 19618 44090 19642 44092
rect 19698 44090 19722 44092
rect 19778 44090 19802 44092
rect 19640 44038 19642 44090
rect 19704 44038 19716 44090
rect 19778 44038 19780 44090
rect 19618 44036 19642 44038
rect 19698 44036 19722 44038
rect 19778 44036 19802 44038
rect 19562 44016 19858 44036
rect 19562 43004 19858 43024
rect 19618 43002 19642 43004
rect 19698 43002 19722 43004
rect 19778 43002 19802 43004
rect 19640 42950 19642 43002
rect 19704 42950 19716 43002
rect 19778 42950 19780 43002
rect 19618 42948 19642 42950
rect 19698 42948 19722 42950
rect 19778 42948 19802 42950
rect 19562 42928 19858 42948
rect 19562 41916 19858 41936
rect 19618 41914 19642 41916
rect 19698 41914 19722 41916
rect 19778 41914 19802 41916
rect 19640 41862 19642 41914
rect 19704 41862 19716 41914
rect 19778 41862 19780 41914
rect 19618 41860 19642 41862
rect 19698 41860 19722 41862
rect 19778 41860 19802 41862
rect 19562 41840 19858 41860
rect 19562 40828 19858 40848
rect 19618 40826 19642 40828
rect 19698 40826 19722 40828
rect 19778 40826 19802 40828
rect 19640 40774 19642 40826
rect 19704 40774 19716 40826
rect 19778 40774 19780 40826
rect 19618 40772 19642 40774
rect 19698 40772 19722 40774
rect 19778 40772 19802 40774
rect 19562 40752 19858 40772
rect 19562 39740 19858 39760
rect 19618 39738 19642 39740
rect 19698 39738 19722 39740
rect 19778 39738 19802 39740
rect 19640 39686 19642 39738
rect 19704 39686 19716 39738
rect 19778 39686 19780 39738
rect 19618 39684 19642 39686
rect 19698 39684 19722 39686
rect 19778 39684 19802 39686
rect 19562 39664 19858 39684
rect 19562 38652 19858 38672
rect 19618 38650 19642 38652
rect 19698 38650 19722 38652
rect 19778 38650 19802 38652
rect 19640 38598 19642 38650
rect 19704 38598 19716 38650
rect 19778 38598 19780 38650
rect 19618 38596 19642 38598
rect 19698 38596 19722 38598
rect 19778 38596 19802 38598
rect 19562 38576 19858 38596
rect 19562 37564 19858 37584
rect 19618 37562 19642 37564
rect 19698 37562 19722 37564
rect 19778 37562 19802 37564
rect 19640 37510 19642 37562
rect 19704 37510 19716 37562
rect 19778 37510 19780 37562
rect 19618 37508 19642 37510
rect 19698 37508 19722 37510
rect 19778 37508 19802 37510
rect 19562 37488 19858 37508
rect 19414 36916 19466 36922
rect 19414 36858 19466 36864
rect 19562 36476 19858 36496
rect 19618 36474 19642 36476
rect 19698 36474 19722 36476
rect 19778 36474 19802 36476
rect 19640 36422 19642 36474
rect 19704 36422 19716 36474
rect 19778 36422 19780 36474
rect 19618 36420 19642 36422
rect 19698 36420 19722 36422
rect 19778 36420 19802 36422
rect 19562 36400 19858 36420
rect 19562 35388 19858 35408
rect 19618 35386 19642 35388
rect 19698 35386 19722 35388
rect 19778 35386 19802 35388
rect 19640 35334 19642 35386
rect 19704 35334 19716 35386
rect 19778 35334 19780 35386
rect 19618 35332 19642 35334
rect 19698 35332 19722 35334
rect 19778 35332 19802 35334
rect 19562 35312 19858 35332
rect 19562 34300 19858 34320
rect 19618 34298 19642 34300
rect 19698 34298 19722 34300
rect 19778 34298 19802 34300
rect 19640 34246 19642 34298
rect 19704 34246 19716 34298
rect 19778 34246 19780 34298
rect 19618 34244 19642 34246
rect 19698 34244 19722 34246
rect 19778 34244 19802 34246
rect 19562 34224 19858 34244
rect 19562 33212 19858 33232
rect 19618 33210 19642 33212
rect 19698 33210 19722 33212
rect 19778 33210 19802 33212
rect 19640 33158 19642 33210
rect 19704 33158 19716 33210
rect 19778 33158 19780 33210
rect 19618 33156 19642 33158
rect 19698 33156 19722 33158
rect 19778 33156 19802 33158
rect 19562 33136 19858 33156
rect 19562 32124 19858 32144
rect 19618 32122 19642 32124
rect 19698 32122 19722 32124
rect 19778 32122 19802 32124
rect 19640 32070 19642 32122
rect 19704 32070 19716 32122
rect 19778 32070 19780 32122
rect 19618 32068 19642 32070
rect 19698 32068 19722 32070
rect 19778 32068 19802 32070
rect 19562 32048 19858 32068
rect 19562 31036 19858 31056
rect 19618 31034 19642 31036
rect 19698 31034 19722 31036
rect 19778 31034 19802 31036
rect 19640 30982 19642 31034
rect 19704 30982 19716 31034
rect 19778 30982 19780 31034
rect 19618 30980 19642 30982
rect 19698 30980 19722 30982
rect 19778 30980 19802 30982
rect 19562 30960 19858 30980
rect 19562 29948 19858 29968
rect 19618 29946 19642 29948
rect 19698 29946 19722 29948
rect 19778 29946 19802 29948
rect 19640 29894 19642 29946
rect 19704 29894 19716 29946
rect 19778 29894 19780 29946
rect 19618 29892 19642 29894
rect 19698 29892 19722 29894
rect 19778 29892 19802 29894
rect 19562 29872 19858 29892
rect 18860 28999 18916 29008
rect 19046 29028 19098 29034
rect 19046 28970 19098 28976
rect 19138 29028 19190 29034
rect 19138 28970 19190 28976
rect 18952 28928 19008 28937
rect 18952 28863 19008 28872
rect 18966 27606 18994 28863
rect 18862 27600 18914 27606
rect 18862 27542 18914 27548
rect 18954 27600 19006 27606
rect 18954 27542 19006 27548
rect 18770 23724 18822 23730
rect 18770 23666 18822 23672
rect 18782 20874 18810 23666
rect 18770 20868 18822 20874
rect 18770 20810 18822 20816
rect 18874 18057 18902 27542
rect 19058 24154 19086 28970
rect 19562 28860 19858 28880
rect 19618 28858 19642 28860
rect 19698 28858 19722 28860
rect 19778 28858 19802 28860
rect 19640 28806 19642 28858
rect 19704 28806 19716 28858
rect 19778 28806 19780 28858
rect 19618 28804 19642 28806
rect 19698 28804 19722 28806
rect 19778 28804 19802 28806
rect 19562 28784 19858 28804
rect 19562 27772 19858 27792
rect 19618 27770 19642 27772
rect 19698 27770 19722 27772
rect 19778 27770 19802 27772
rect 19640 27718 19642 27770
rect 19704 27718 19716 27770
rect 19778 27718 19780 27770
rect 19618 27716 19642 27718
rect 19698 27716 19722 27718
rect 19778 27716 19802 27718
rect 19562 27696 19858 27716
rect 19562 26684 19858 26704
rect 19618 26682 19642 26684
rect 19698 26682 19722 26684
rect 19778 26682 19802 26684
rect 19640 26630 19642 26682
rect 19704 26630 19716 26682
rect 19778 26630 19780 26682
rect 19618 26628 19642 26630
rect 19698 26628 19722 26630
rect 19778 26628 19802 26630
rect 19562 26608 19858 26628
rect 19562 25596 19858 25616
rect 19618 25594 19642 25596
rect 19698 25594 19722 25596
rect 19778 25594 19802 25596
rect 19640 25542 19642 25594
rect 19704 25542 19716 25594
rect 19778 25542 19780 25594
rect 19618 25540 19642 25542
rect 19698 25540 19722 25542
rect 19778 25540 19802 25542
rect 19562 25520 19858 25540
rect 19562 24508 19858 24528
rect 19618 24506 19642 24508
rect 19698 24506 19722 24508
rect 19778 24506 19802 24508
rect 19640 24454 19642 24506
rect 19704 24454 19716 24506
rect 19778 24454 19780 24506
rect 19618 24452 19642 24454
rect 19698 24452 19722 24454
rect 19778 24452 19802 24454
rect 19562 24432 19858 24452
rect 19058 24126 19270 24154
rect 18860 18048 18916 18057
rect 18860 17983 18916 17992
rect 18952 17912 19008 17921
rect 18952 17847 19008 17856
rect 18678 15088 18730 15094
rect 18678 15030 18730 15036
rect 18862 14544 18914 14550
rect 18862 14486 18914 14492
rect 18770 7540 18822 7546
rect 18770 7482 18822 7488
rect 18586 3188 18638 3194
rect 18586 3130 18638 3136
rect 18586 3052 18638 3058
rect 18586 2994 18638 3000
rect 18598 800 18626 2994
rect 18782 800 18810 7482
rect 18874 4146 18902 14486
rect 18966 6322 18994 17847
rect 19046 11688 19098 11694
rect 19046 11630 19098 11636
rect 18954 6316 19006 6322
rect 18954 6258 19006 6264
rect 18954 4208 19006 4214
rect 18954 4150 19006 4156
rect 18862 4140 18914 4146
rect 18862 4082 18914 4088
rect 18966 3777 18994 4150
rect 18952 3768 19008 3777
rect 18952 3703 19008 3712
rect 19058 3126 19086 11630
rect 19242 3890 19270 24126
rect 19562 23420 19858 23440
rect 19618 23418 19642 23420
rect 19698 23418 19722 23420
rect 19778 23418 19802 23420
rect 19640 23366 19642 23418
rect 19704 23366 19716 23418
rect 19778 23366 19780 23418
rect 19618 23364 19642 23366
rect 19698 23364 19722 23366
rect 19778 23364 19802 23366
rect 19562 23344 19858 23364
rect 19562 22332 19858 22352
rect 19618 22330 19642 22332
rect 19698 22330 19722 22332
rect 19778 22330 19802 22332
rect 19640 22278 19642 22330
rect 19704 22278 19716 22330
rect 19778 22278 19780 22330
rect 19618 22276 19642 22278
rect 19698 22276 19722 22278
rect 19778 22276 19802 22278
rect 19562 22256 19858 22276
rect 19562 21244 19858 21264
rect 19618 21242 19642 21244
rect 19698 21242 19722 21244
rect 19778 21242 19802 21244
rect 19640 21190 19642 21242
rect 19704 21190 19716 21242
rect 19778 21190 19780 21242
rect 19618 21188 19642 21190
rect 19698 21188 19722 21190
rect 19778 21188 19802 21190
rect 19562 21168 19858 21188
rect 19562 20156 19858 20176
rect 19618 20154 19642 20156
rect 19698 20154 19722 20156
rect 19778 20154 19802 20156
rect 19640 20102 19642 20154
rect 19704 20102 19716 20154
rect 19778 20102 19780 20154
rect 19618 20100 19642 20102
rect 19698 20100 19722 20102
rect 19778 20100 19802 20102
rect 19562 20080 19858 20100
rect 19562 19068 19858 19088
rect 19618 19066 19642 19068
rect 19698 19066 19722 19068
rect 19778 19066 19802 19068
rect 19640 19014 19642 19066
rect 19704 19014 19716 19066
rect 19778 19014 19780 19066
rect 19618 19012 19642 19014
rect 19698 19012 19722 19014
rect 19778 19012 19802 19014
rect 19562 18992 19858 19012
rect 19562 17980 19858 18000
rect 19618 17978 19642 17980
rect 19698 17978 19722 17980
rect 19778 17978 19802 17980
rect 19640 17926 19642 17978
rect 19704 17926 19716 17978
rect 19778 17926 19780 17978
rect 19618 17924 19642 17926
rect 19698 17924 19722 17926
rect 19778 17924 19802 17926
rect 19562 17904 19858 17924
rect 19322 17536 19374 17542
rect 19320 17504 19322 17513
rect 19374 17504 19376 17513
rect 19320 17439 19376 17448
rect 19562 16892 19858 16912
rect 19618 16890 19642 16892
rect 19698 16890 19722 16892
rect 19778 16890 19802 16892
rect 19640 16838 19642 16890
rect 19704 16838 19716 16890
rect 19778 16838 19780 16890
rect 19618 16836 19642 16838
rect 19698 16836 19722 16838
rect 19778 16836 19802 16838
rect 19562 16816 19858 16836
rect 19562 15804 19858 15824
rect 19618 15802 19642 15804
rect 19698 15802 19722 15804
rect 19778 15802 19802 15804
rect 19640 15750 19642 15802
rect 19704 15750 19716 15802
rect 19778 15750 19780 15802
rect 19618 15748 19642 15750
rect 19698 15748 19722 15750
rect 19778 15748 19802 15750
rect 19562 15728 19858 15748
rect 19562 14716 19858 14736
rect 19618 14714 19642 14716
rect 19698 14714 19722 14716
rect 19778 14714 19802 14716
rect 19640 14662 19642 14714
rect 19704 14662 19716 14714
rect 19778 14662 19780 14714
rect 19618 14660 19642 14662
rect 19698 14660 19722 14662
rect 19778 14660 19802 14662
rect 19562 14640 19858 14660
rect 19562 13628 19858 13648
rect 19618 13626 19642 13628
rect 19698 13626 19722 13628
rect 19778 13626 19802 13628
rect 19640 13574 19642 13626
rect 19704 13574 19716 13626
rect 19778 13574 19780 13626
rect 19618 13572 19642 13574
rect 19698 13572 19722 13574
rect 19778 13572 19802 13574
rect 19562 13552 19858 13572
rect 19562 12540 19858 12560
rect 19618 12538 19642 12540
rect 19698 12538 19722 12540
rect 19778 12538 19802 12540
rect 19640 12486 19642 12538
rect 19704 12486 19716 12538
rect 19778 12486 19780 12538
rect 19618 12484 19642 12486
rect 19698 12484 19722 12486
rect 19778 12484 19802 12486
rect 19562 12464 19858 12484
rect 19562 11452 19858 11472
rect 19618 11450 19642 11452
rect 19698 11450 19722 11452
rect 19778 11450 19802 11452
rect 19640 11398 19642 11450
rect 19704 11398 19716 11450
rect 19778 11398 19780 11450
rect 19618 11396 19642 11398
rect 19698 11396 19722 11398
rect 19778 11396 19802 11398
rect 19562 11376 19858 11396
rect 19562 10364 19858 10384
rect 19618 10362 19642 10364
rect 19698 10362 19722 10364
rect 19778 10362 19802 10364
rect 19640 10310 19642 10362
rect 19704 10310 19716 10362
rect 19778 10310 19780 10362
rect 19618 10308 19642 10310
rect 19698 10308 19722 10310
rect 19778 10308 19802 10310
rect 19562 10288 19858 10308
rect 19562 9276 19858 9296
rect 19618 9274 19642 9276
rect 19698 9274 19722 9276
rect 19778 9274 19802 9276
rect 19640 9222 19642 9274
rect 19704 9222 19716 9274
rect 19778 9222 19780 9274
rect 19618 9220 19642 9222
rect 19698 9220 19722 9222
rect 19778 9220 19802 9222
rect 19562 9200 19858 9220
rect 19562 8188 19858 8208
rect 19618 8186 19642 8188
rect 19698 8186 19722 8188
rect 19778 8186 19802 8188
rect 19640 8134 19642 8186
rect 19704 8134 19716 8186
rect 19778 8134 19780 8186
rect 19618 8132 19642 8134
rect 19698 8132 19722 8134
rect 19778 8132 19802 8134
rect 19562 8112 19858 8132
rect 19886 7721 19914 53638
rect 20070 53122 20098 55286
rect 19978 53094 20098 53122
rect 19978 41274 20006 53094
rect 20058 43648 20110 43654
rect 20058 43590 20110 43596
rect 19966 41268 20018 41274
rect 19966 41210 20018 41216
rect 19966 20868 20018 20874
rect 19966 20810 20018 20816
rect 19872 7712 19928 7721
rect 19872 7647 19928 7656
rect 19872 7576 19928 7585
rect 19414 7540 19466 7546
rect 19872 7511 19928 7520
rect 19414 7482 19466 7488
rect 19322 4140 19374 4146
rect 19322 4082 19374 4088
rect 19150 3862 19270 3890
rect 19046 3120 19098 3126
rect 19046 3062 19098 3068
rect 19150 2938 19178 3862
rect 18966 2910 19178 2938
rect 18966 800 18994 2910
rect 19334 800 19362 4082
rect 19426 1442 19454 7482
rect 19562 7100 19858 7120
rect 19618 7098 19642 7100
rect 19698 7098 19722 7100
rect 19778 7098 19802 7100
rect 19640 7046 19642 7098
rect 19704 7046 19716 7098
rect 19778 7046 19780 7098
rect 19618 7044 19642 7046
rect 19698 7044 19722 7046
rect 19778 7044 19802 7046
rect 19562 7024 19858 7044
rect 19562 6012 19858 6032
rect 19618 6010 19642 6012
rect 19698 6010 19722 6012
rect 19778 6010 19802 6012
rect 19640 5958 19642 6010
rect 19704 5958 19716 6010
rect 19778 5958 19780 6010
rect 19618 5956 19642 5958
rect 19698 5956 19722 5958
rect 19778 5956 19802 5958
rect 19562 5936 19858 5956
rect 19562 4924 19858 4944
rect 19618 4922 19642 4924
rect 19698 4922 19722 4924
rect 19778 4922 19802 4924
rect 19640 4870 19642 4922
rect 19704 4870 19716 4922
rect 19778 4870 19780 4922
rect 19618 4868 19642 4870
rect 19698 4868 19722 4870
rect 19778 4868 19802 4870
rect 19562 4848 19858 4868
rect 19562 3836 19858 3856
rect 19618 3834 19642 3836
rect 19698 3834 19722 3836
rect 19778 3834 19802 3836
rect 19640 3782 19642 3834
rect 19704 3782 19716 3834
rect 19778 3782 19780 3834
rect 19618 3780 19642 3782
rect 19698 3780 19722 3782
rect 19778 3780 19802 3782
rect 19562 3760 19858 3780
rect 19562 2748 19858 2768
rect 19618 2746 19642 2748
rect 19698 2746 19722 2748
rect 19778 2746 19802 2748
rect 19640 2694 19642 2746
rect 19704 2694 19716 2746
rect 19778 2694 19780 2746
rect 19618 2692 19642 2694
rect 19698 2692 19722 2694
rect 19778 2692 19802 2694
rect 19562 2672 19858 2692
rect 19426 1414 19546 1442
rect 19518 800 19546 1414
rect 19690 1420 19742 1426
rect 19690 1362 19742 1368
rect 19702 800 19730 1362
rect 19886 800 19914 7511
rect 19978 4078 20006 20810
rect 20070 7426 20098 43590
rect 20162 43178 20190 55762
rect 20530 46510 20558 55950
rect 20714 55418 20742 59200
rect 21070 56432 21122 56438
rect 21070 56374 21122 56380
rect 21082 55622 21110 56374
rect 20978 55616 21030 55622
rect 20978 55558 21030 55564
rect 21070 55616 21122 55622
rect 21070 55558 21122 55564
rect 20702 55412 20754 55418
rect 20702 55354 20754 55360
rect 20990 55350 21018 55558
rect 20978 55344 21030 55350
rect 20978 55286 21030 55292
rect 20610 55276 20662 55282
rect 20610 55218 20662 55224
rect 20518 46504 20570 46510
rect 20518 46446 20570 46452
rect 20518 45824 20570 45830
rect 20518 45766 20570 45772
rect 20530 45626 20558 45766
rect 20518 45620 20570 45626
rect 20518 45562 20570 45568
rect 20150 43172 20202 43178
rect 20150 43114 20202 43120
rect 20518 39432 20570 39438
rect 20518 39374 20570 39380
rect 20334 25900 20386 25906
rect 20334 25842 20386 25848
rect 20346 25770 20374 25842
rect 20334 25764 20386 25770
rect 20334 25706 20386 25712
rect 20426 25764 20478 25770
rect 20426 25706 20478 25712
rect 20334 24132 20386 24138
rect 20334 24074 20386 24080
rect 20150 23656 20202 23662
rect 20150 23598 20202 23604
rect 20162 7585 20190 23598
rect 20242 23520 20294 23526
rect 20242 23462 20294 23468
rect 20148 7576 20204 7585
rect 20148 7511 20204 7520
rect 20070 7398 20190 7426
rect 20058 4140 20110 4146
rect 20058 4082 20110 4088
rect 19966 4072 20018 4078
rect 19966 4014 20018 4020
rect 20070 800 20098 4082
rect 20162 4010 20190 7398
rect 20150 4004 20202 4010
rect 20150 3946 20202 3952
rect 20254 800 20282 23462
rect 20346 7546 20374 24074
rect 20334 7540 20386 7546
rect 20334 7482 20386 7488
rect 20438 4146 20466 25706
rect 20426 4140 20478 4146
rect 20426 4082 20478 4088
rect 20530 1426 20558 39374
rect 20622 5914 20650 55218
rect 21174 52034 21202 59200
rect 21622 56228 21674 56234
rect 21622 56170 21674 56176
rect 21634 53666 21662 56170
rect 21726 54262 21754 59200
rect 22738 55690 22766 59200
rect 22726 55684 22778 55690
rect 22726 55626 22778 55632
rect 23290 55622 23318 59200
rect 23738 56840 23790 56846
rect 23738 56782 23790 56788
rect 23750 56506 23778 56782
rect 23738 56500 23790 56506
rect 23738 56442 23790 56448
rect 23278 55616 23330 55622
rect 23278 55558 23330 55564
rect 23370 55412 23422 55418
rect 23370 55354 23422 55360
rect 22542 54528 22594 54534
rect 22542 54470 22594 54476
rect 22554 54330 22582 54470
rect 22542 54324 22594 54330
rect 22542 54266 22594 54272
rect 21714 54256 21766 54262
rect 21714 54198 21766 54204
rect 22726 54120 22778 54126
rect 22726 54062 22778 54068
rect 21634 53638 21846 53666
rect 21082 52006 21202 52034
rect 20702 26920 20754 26926
rect 20702 26862 20754 26868
rect 20714 19242 20742 26862
rect 20886 24812 20938 24818
rect 20886 24754 20938 24760
rect 20702 19236 20754 19242
rect 20702 19178 20754 19184
rect 20702 8424 20754 8430
rect 20702 8366 20754 8372
rect 20610 5908 20662 5914
rect 20610 5850 20662 5856
rect 20714 2990 20742 8366
rect 20898 4842 20926 24754
rect 20978 24744 21030 24750
rect 20978 24686 21030 24692
rect 20990 5030 21018 24686
rect 21082 12442 21110 52006
rect 21346 45892 21398 45898
rect 21346 45834 21398 45840
rect 21358 19446 21386 45834
rect 21818 37466 21846 53638
rect 21806 37460 21858 37466
rect 21806 37402 21858 37408
rect 21438 35624 21490 35630
rect 21438 35566 21490 35572
rect 21346 19440 21398 19446
rect 21346 19382 21398 19388
rect 21162 19304 21214 19310
rect 21162 19246 21214 19252
rect 21070 12436 21122 12442
rect 21070 12378 21122 12384
rect 21070 8084 21122 8090
rect 21070 8026 21122 8032
rect 20978 5024 21030 5030
rect 20978 4966 21030 4972
rect 20898 4814 21018 4842
rect 20794 4072 20846 4078
rect 20794 4014 20846 4020
rect 20702 2984 20754 2990
rect 20702 2926 20754 2932
rect 20518 1420 20570 1426
rect 20518 1362 20570 1368
rect 20424 912 20480 921
rect 20424 847 20480 856
rect 20438 800 20466 847
rect 20806 800 20834 4014
rect 20990 2802 21018 4814
rect 21082 3058 21110 8026
rect 21174 4282 21202 19246
rect 21346 12844 21398 12850
rect 21346 12786 21398 12792
rect 21358 12714 21386 12786
rect 21346 12708 21398 12714
rect 21346 12650 21398 12656
rect 21346 10124 21398 10130
rect 21346 10066 21398 10072
rect 21358 9926 21386 10066
rect 21346 9920 21398 9926
rect 21346 9862 21398 9868
rect 21450 8430 21478 35566
rect 22634 32972 22686 32978
rect 22634 32914 22686 32920
rect 22646 32774 22674 32914
rect 22634 32768 22686 32774
rect 22634 32710 22686 32716
rect 21990 31816 22042 31822
rect 21990 31758 22042 31764
rect 21622 25424 21674 25430
rect 21622 25366 21674 25372
rect 21530 24948 21582 24954
rect 21530 24890 21582 24896
rect 21438 8424 21490 8430
rect 21438 8366 21490 8372
rect 21542 8242 21570 24890
rect 21266 8214 21570 8242
rect 21162 4276 21214 4282
rect 21162 4218 21214 4224
rect 21266 4146 21294 8214
rect 21634 8090 21662 25366
rect 21714 24676 21766 24682
rect 21714 24618 21766 24624
rect 21622 8084 21674 8090
rect 21622 8026 21674 8032
rect 21726 7970 21754 24618
rect 21806 24404 21858 24410
rect 21806 24346 21858 24352
rect 21450 7942 21754 7970
rect 21346 7744 21398 7750
rect 21346 7686 21398 7692
rect 21254 4140 21306 4146
rect 21254 4082 21306 4088
rect 21162 4004 21214 4010
rect 21162 3946 21214 3952
rect 21254 4004 21306 4010
rect 21254 3946 21306 3952
rect 21070 3052 21122 3058
rect 21070 2994 21122 3000
rect 20990 2774 21110 2802
rect 21082 898 21110 2774
rect 20990 870 21110 898
rect 20990 800 21018 870
rect 21174 800 21202 3946
rect 21266 3398 21294 3946
rect 21254 3392 21306 3398
rect 21254 3334 21306 3340
rect 21358 800 21386 7686
rect 21450 3398 21478 7942
rect 21818 7750 21846 24346
rect 21898 12844 21950 12850
rect 21898 12786 21950 12792
rect 21806 7744 21858 7750
rect 21806 7686 21858 7692
rect 21910 7562 21938 12786
rect 21542 7534 21938 7562
rect 21438 3392 21490 3398
rect 21438 3334 21490 3340
rect 21542 800 21570 7534
rect 21714 5024 21766 5030
rect 21714 4966 21766 4972
rect 21726 800 21754 4966
rect 22002 4842 22030 31758
rect 22450 25696 22502 25702
rect 22450 25638 22502 25644
rect 22358 7880 22410 7886
rect 22358 7822 22410 7828
rect 21818 4814 22030 4842
rect 21818 2666 21846 4814
rect 22266 4276 22318 4282
rect 22266 4218 22318 4224
rect 22082 3392 22134 3398
rect 22082 3334 22134 3340
rect 21818 2638 21938 2666
rect 21910 800 21938 2638
rect 22094 800 22122 3334
rect 22278 800 22306 4218
rect 22370 2922 22398 7822
rect 22358 2916 22410 2922
rect 22358 2858 22410 2864
rect 22462 2650 22490 25638
rect 22634 25492 22686 25498
rect 22634 25434 22686 25440
rect 22646 7750 22674 25434
rect 22738 7886 22766 54062
rect 23382 53242 23410 55354
rect 23842 55162 23870 59200
rect 24014 56296 24066 56302
rect 24014 56238 24066 56244
rect 24026 55350 24054 56238
rect 24014 55344 24066 55350
rect 24014 55286 24066 55292
rect 23474 55134 23870 55162
rect 24394 55162 24422 59200
rect 24854 55282 24882 59200
rect 25958 55622 25986 59200
rect 26038 56704 26090 56710
rect 26038 56646 26090 56652
rect 25946 55616 25998 55622
rect 25946 55558 25998 55564
rect 26050 55400 26078 56646
rect 26222 55820 26274 55826
rect 26222 55762 26274 55768
rect 26234 55690 26262 55762
rect 26222 55684 26274 55690
rect 26222 55626 26274 55632
rect 25958 55372 26078 55400
rect 24842 55276 24894 55282
rect 24842 55218 24894 55224
rect 24394 55134 24790 55162
rect 23370 53236 23422 53242
rect 23370 53178 23422 53184
rect 23186 45824 23238 45830
rect 23186 45766 23238 45772
rect 23198 44169 23226 45766
rect 23000 44160 23056 44169
rect 23000 44095 23056 44104
rect 23184 44160 23240 44169
rect 23184 44095 23240 44104
rect 23014 34542 23042 44095
rect 23370 43648 23422 43654
rect 23370 43590 23422 43596
rect 23382 39438 23410 43590
rect 23370 39432 23422 39438
rect 23370 39374 23422 39380
rect 23002 34536 23054 34542
rect 23002 34478 23054 34484
rect 23186 34536 23238 34542
rect 23186 34478 23238 34484
rect 23198 32502 23226 34478
rect 23186 32496 23238 32502
rect 23186 32438 23238 32444
rect 23474 28694 23502 55134
rect 23552 54632 23608 54641
rect 23552 54567 23608 54576
rect 23566 54534 23594 54567
rect 23554 54528 23606 54534
rect 23554 54470 23606 54476
rect 24198 48340 24250 48346
rect 24198 48282 24250 48288
rect 24210 41154 24238 48282
rect 24118 41126 24238 41154
rect 24118 38729 24146 41126
rect 24198 40996 24250 41002
rect 24198 40938 24250 40944
rect 24104 38720 24160 38729
rect 24104 38655 24160 38664
rect 24104 38584 24160 38593
rect 24104 38519 24160 38528
rect 23554 32496 23606 32502
rect 23554 32438 23606 32444
rect 23278 28688 23330 28694
rect 23278 28630 23330 28636
rect 23462 28688 23514 28694
rect 23462 28630 23514 28636
rect 22818 27872 22870 27878
rect 22818 27814 22870 27820
rect 22830 7954 22858 27814
rect 23002 26852 23054 26858
rect 23002 26794 23054 26800
rect 22910 26580 22962 26586
rect 22910 26522 22962 26528
rect 22818 7948 22870 7954
rect 22818 7890 22870 7896
rect 22726 7880 22778 7886
rect 22922 7834 22950 26522
rect 22726 7822 22778 7828
rect 22830 7806 22950 7834
rect 22634 7744 22686 7750
rect 22634 7686 22686 7692
rect 22634 4140 22686 4146
rect 22634 4082 22686 4088
rect 22542 4004 22594 4010
rect 22542 3946 22594 3952
rect 22554 3194 22582 3946
rect 22542 3188 22594 3194
rect 22542 3130 22594 3136
rect 22450 2644 22502 2650
rect 22450 2586 22502 2592
rect 22646 800 22674 4082
rect 22830 4078 22858 7806
rect 22910 7744 22962 7750
rect 22910 7686 22962 7692
rect 23014 7698 23042 26794
rect 23290 24954 23318 28630
rect 23278 24948 23330 24954
rect 23278 24890 23330 24896
rect 23462 24948 23514 24954
rect 23462 24890 23514 24896
rect 23186 19236 23238 19242
rect 23186 19178 23238 19184
rect 22818 4072 22870 4078
rect 22818 4014 22870 4020
rect 22922 2650 22950 7686
rect 23014 7670 23134 7698
rect 23002 7540 23054 7546
rect 23002 7482 23054 7488
rect 22818 2644 22870 2650
rect 22818 2586 22870 2592
rect 22910 2644 22962 2650
rect 22910 2586 22962 2592
rect 22830 800 22858 2586
rect 23014 800 23042 7482
rect 23106 3398 23134 7670
rect 23198 3738 23226 19178
rect 23370 17332 23422 17338
rect 23370 17274 23422 17280
rect 23382 17241 23410 17274
rect 23368 17232 23424 17241
rect 23368 17167 23424 17176
rect 23276 15192 23332 15201
rect 23276 15127 23332 15136
rect 23290 7546 23318 15127
rect 23370 7948 23422 7954
rect 23370 7890 23422 7896
rect 23278 7540 23330 7546
rect 23278 7482 23330 7488
rect 23186 3732 23238 3738
rect 23186 3674 23238 3680
rect 23094 3392 23146 3398
rect 23094 3334 23146 3340
rect 23382 3126 23410 7890
rect 23474 7410 23502 24890
rect 23566 23361 23594 32438
rect 24118 29034 24146 38519
rect 24014 29028 24066 29034
rect 24014 28970 24066 28976
rect 24106 29028 24158 29034
rect 24106 28970 24158 28976
rect 23552 23352 23608 23361
rect 23552 23287 23608 23296
rect 24026 22794 24054 28970
rect 24026 22766 24146 22794
rect 23830 12776 23882 12782
rect 23830 12718 23882 12724
rect 23462 7404 23514 7410
rect 23462 7346 23514 7352
rect 23842 4554 23870 12718
rect 24014 10124 24066 10130
rect 24014 10066 24066 10072
rect 24026 9994 24054 10066
rect 24014 9988 24066 9994
rect 24014 9930 24066 9936
rect 24014 8628 24066 8634
rect 24014 8570 24066 8576
rect 23830 4548 23882 4554
rect 23830 4490 23882 4496
rect 23922 3392 23974 3398
rect 23922 3334 23974 3340
rect 23370 3120 23422 3126
rect 23370 3062 23422 3068
rect 23738 3052 23790 3058
rect 23738 2994 23790 3000
rect 23370 2984 23422 2990
rect 23370 2926 23422 2932
rect 23186 2644 23238 2650
rect 23186 2586 23238 2592
rect 23198 800 23226 2586
rect 23382 800 23410 2926
rect 23750 800 23778 2994
rect 23934 800 23962 3334
rect 24026 2836 24054 8570
rect 24118 7206 24146 22766
rect 24106 7200 24158 7206
rect 24106 7142 24158 7148
rect 24210 3058 24238 40938
rect 24382 28960 24434 28966
rect 24382 28902 24434 28908
rect 24290 28008 24342 28014
rect 24290 27950 24342 27956
rect 24302 4146 24330 27950
rect 24290 4140 24342 4146
rect 24290 4082 24342 4088
rect 24290 3732 24342 3738
rect 24290 3674 24342 3680
rect 24198 3052 24250 3058
rect 24198 2994 24250 3000
rect 24026 2808 24146 2836
rect 24118 800 24146 2808
rect 24302 800 24330 3674
rect 24394 3398 24422 28902
rect 24658 26852 24710 26858
rect 24658 26794 24710 26800
rect 24566 17536 24618 17542
rect 24564 17504 24566 17513
rect 24618 17504 24620 17513
rect 24564 17439 24620 17448
rect 24566 17128 24618 17134
rect 24566 17070 24618 17076
rect 24578 16114 24606 17070
rect 24566 16108 24618 16114
rect 24566 16050 24618 16056
rect 24670 4842 24698 26794
rect 24762 17134 24790 55134
rect 25958 46170 25986 55372
rect 26038 55276 26090 55282
rect 26038 55218 26090 55224
rect 25946 46164 25998 46170
rect 25946 46106 25998 46112
rect 25946 36372 25998 36378
rect 25946 36314 25998 36320
rect 25486 30048 25538 30054
rect 25486 29990 25538 29996
rect 25394 28076 25446 28082
rect 25394 28018 25446 28024
rect 25026 26308 25078 26314
rect 25026 26250 25078 26256
rect 24750 17128 24802 17134
rect 24750 17070 24802 17076
rect 24934 16176 24986 16182
rect 24934 16118 24986 16124
rect 24946 15978 24974 16118
rect 24750 15972 24802 15978
rect 24750 15914 24802 15920
rect 24934 15972 24986 15978
rect 24934 15914 24986 15920
rect 24762 15881 24790 15914
rect 24748 15872 24804 15881
rect 24748 15807 24804 15816
rect 24748 11656 24804 11665
rect 24804 11626 24882 11642
rect 24804 11620 24894 11626
rect 24804 11614 24842 11620
rect 24748 11591 24804 11600
rect 24842 11562 24894 11568
rect 24842 10804 24894 10810
rect 24842 10746 24894 10752
rect 24854 10690 24882 10746
rect 24762 10662 24882 10690
rect 24762 10606 24790 10662
rect 24750 10600 24802 10606
rect 24750 10542 24802 10548
rect 24486 4814 24698 4842
rect 24382 3392 24434 3398
rect 24382 3334 24434 3340
rect 24486 800 24514 4814
rect 25038 4282 25066 26250
rect 25118 7744 25170 7750
rect 25118 7686 25170 7692
rect 25130 7478 25158 7686
rect 25118 7472 25170 7478
rect 25118 7414 25170 7420
rect 25026 4276 25078 4282
rect 25026 4218 25078 4224
rect 25026 4140 25078 4146
rect 25026 4082 25078 4088
rect 25210 4140 25262 4146
rect 25210 4082 25262 4088
rect 24842 4072 24894 4078
rect 24842 4014 24894 4020
rect 24854 800 24882 4014
rect 25038 800 25066 4082
rect 25222 800 25250 4082
rect 25406 800 25434 28018
rect 25498 4010 25526 29990
rect 25854 29572 25906 29578
rect 25854 29514 25906 29520
rect 25670 14408 25722 14414
rect 25670 14350 25722 14356
rect 25578 7744 25630 7750
rect 25578 7686 25630 7692
rect 25486 4004 25538 4010
rect 25486 3946 25538 3952
rect 25590 800 25618 7686
rect 25682 2650 25710 14350
rect 25762 14272 25814 14278
rect 25762 14214 25814 14220
rect 25774 14074 25802 14214
rect 25762 14068 25814 14074
rect 25762 14010 25814 14016
rect 25866 4026 25894 29514
rect 25958 26926 25986 36314
rect 25946 26920 25998 26926
rect 25946 26862 25998 26868
rect 25946 22568 25998 22574
rect 25946 22510 25998 22516
rect 25958 7750 25986 22510
rect 26050 19718 26078 55218
rect 26418 48346 26446 59200
rect 26970 56817 26998 59200
rect 26956 56808 27012 56817
rect 26956 56743 27012 56752
rect 26864 56672 26920 56681
rect 26920 56630 26998 56658
rect 26864 56607 26920 56616
rect 26680 56400 26736 56409
rect 26680 56335 26682 56344
rect 26734 56335 26736 56344
rect 26774 56364 26826 56370
rect 26682 56306 26734 56312
rect 26774 56306 26826 56312
rect 26786 55758 26814 56306
rect 26866 56228 26918 56234
rect 26866 56170 26918 56176
rect 26878 55758 26906 56170
rect 26774 55752 26826 55758
rect 26774 55694 26826 55700
rect 26866 55752 26918 55758
rect 26866 55694 26918 55700
rect 26970 48362 26998 56630
rect 27050 56228 27102 56234
rect 27050 56170 27102 56176
rect 26406 48340 26458 48346
rect 26406 48282 26458 48288
rect 26878 48334 26998 48362
rect 26878 47054 26906 48334
rect 26866 47048 26918 47054
rect 26866 46990 26918 46996
rect 26590 46980 26642 46986
rect 26590 46922 26642 46928
rect 26130 46164 26182 46170
rect 26130 46106 26182 46112
rect 26142 36378 26170 46106
rect 26602 45558 26630 46922
rect 26222 45552 26274 45558
rect 26222 45494 26274 45500
rect 26590 45552 26642 45558
rect 26590 45494 26642 45500
rect 26130 36372 26182 36378
rect 26130 36314 26182 36320
rect 26234 36038 26262 45494
rect 26866 44396 26918 44402
rect 26866 44338 26918 44344
rect 26222 36032 26274 36038
rect 26222 35974 26274 35980
rect 26406 36032 26458 36038
rect 26406 35974 26458 35980
rect 26314 29164 26366 29170
rect 26314 29106 26366 29112
rect 26130 26920 26182 26926
rect 26130 26862 26182 26868
rect 26038 19712 26090 19718
rect 26038 19654 26090 19660
rect 25946 7744 25998 7750
rect 25946 7686 25998 7692
rect 26142 4146 26170 26862
rect 26326 22794 26354 29106
rect 26418 27674 26446 35974
rect 26406 27668 26458 27674
rect 26406 27610 26458 27616
rect 26498 27668 26550 27674
rect 26498 27610 26550 27616
rect 26510 22982 26538 27610
rect 26498 22976 26550 22982
rect 26498 22918 26550 22924
rect 26682 22976 26734 22982
rect 26682 22918 26734 22924
rect 26326 22766 26538 22794
rect 26222 12300 26274 12306
rect 26222 12242 26274 12248
rect 26234 12170 26262 12242
rect 26222 12164 26274 12170
rect 26222 12106 26274 12112
rect 26222 11756 26274 11762
rect 26222 11698 26274 11704
rect 26234 11626 26262 11698
rect 26222 11620 26274 11626
rect 26222 11562 26274 11568
rect 26222 10804 26274 10810
rect 26222 10746 26274 10752
rect 26234 10674 26262 10746
rect 26222 10668 26274 10674
rect 26222 10610 26274 10616
rect 26222 6180 26274 6186
rect 26222 6122 26274 6128
rect 26130 4140 26182 4146
rect 26130 4082 26182 4088
rect 25866 3998 26170 4026
rect 25946 3120 25998 3126
rect 25946 3062 25998 3068
rect 25670 2644 25722 2650
rect 25670 2586 25722 2592
rect 25958 800 25986 3062
rect 26142 800 26170 3998
rect 26234 2990 26262 6122
rect 26314 4140 26366 4146
rect 26314 4082 26366 4088
rect 26222 2984 26274 2990
rect 26222 2926 26274 2932
rect 26326 800 26354 4082
rect 26510 800 26538 22766
rect 26694 8650 26722 22918
rect 26602 8622 26722 8650
rect 26602 8498 26630 8622
rect 26590 8492 26642 8498
rect 26590 8434 26642 8440
rect 26878 7562 26906 44338
rect 26958 32428 27010 32434
rect 26958 32370 27010 32376
rect 26970 19378 26998 32370
rect 27062 23866 27090 56170
rect 27522 55690 27550 59200
rect 28074 56438 28102 59200
rect 28062 56432 28114 56438
rect 28154 56432 28206 56438
rect 28062 56374 28114 56380
rect 28152 56400 28154 56409
rect 28206 56400 28208 56409
rect 28152 56335 28208 56344
rect 27510 55684 27562 55690
rect 27510 55626 27562 55632
rect 27418 55616 27470 55622
rect 27416 55584 27418 55593
rect 27602 55616 27654 55622
rect 27470 55584 27472 55593
rect 27602 55558 27654 55564
rect 27416 55519 27472 55528
rect 27142 54256 27194 54262
rect 27142 54198 27194 54204
rect 27154 46986 27182 54198
rect 27142 46980 27194 46986
rect 27142 46922 27194 46928
rect 27142 40384 27194 40390
rect 27142 40326 27194 40332
rect 27154 32434 27182 40326
rect 27510 39432 27562 39438
rect 27510 39374 27562 39380
rect 27142 32428 27194 32434
rect 27142 32370 27194 32376
rect 27234 29844 27286 29850
rect 27234 29786 27286 29792
rect 27142 29300 27194 29306
rect 27142 29242 27194 29248
rect 27050 23860 27102 23866
rect 27050 23802 27102 23808
rect 26958 19372 27010 19378
rect 26958 19314 27010 19320
rect 27050 19304 27102 19310
rect 27050 19246 27102 19252
rect 26958 8628 27010 8634
rect 26958 8570 27010 8576
rect 26970 8498 26998 8570
rect 26958 8492 27010 8498
rect 26958 8434 27010 8440
rect 26878 7534 26998 7562
rect 26864 3360 26920 3369
rect 26864 3295 26920 3304
rect 26682 2916 26734 2922
rect 26682 2858 26734 2864
rect 26694 800 26722 2858
rect 26878 2825 26906 3295
rect 26970 3126 26998 7534
rect 27062 4078 27090 19246
rect 27050 4072 27102 4078
rect 27050 4014 27102 4020
rect 27050 3392 27102 3398
rect 27050 3334 27102 3340
rect 26958 3120 27010 3126
rect 26958 3062 27010 3068
rect 26864 2816 26920 2825
rect 26864 2751 26920 2760
rect 27062 800 27090 3334
rect 27154 2854 27182 29242
rect 27142 2848 27194 2854
rect 27142 2790 27194 2796
rect 27246 800 27274 29786
rect 27326 19848 27378 19854
rect 27378 19796 27458 19802
rect 27326 19790 27458 19796
rect 27338 19774 27458 19790
rect 27430 19718 27458 19774
rect 27418 19712 27470 19718
rect 27418 19654 27470 19660
rect 27418 4208 27470 4214
rect 27418 4150 27470 4156
rect 27430 3720 27458 4150
rect 27522 4146 27550 39374
rect 27614 28762 27642 55558
rect 29086 55350 29114 59200
rect 29442 56840 29494 56846
rect 29442 56782 29494 56788
rect 29454 56302 29482 56782
rect 29442 56296 29494 56302
rect 29442 56238 29494 56244
rect 29074 55344 29126 55350
rect 29074 55286 29126 55292
rect 29638 55282 29666 59200
rect 29718 56296 29770 56302
rect 29718 56238 29770 56244
rect 28246 55276 28298 55282
rect 28246 55218 28298 55224
rect 29626 55276 29678 55282
rect 29626 55218 29678 55224
rect 27878 30932 27930 30938
rect 27878 30874 27930 30880
rect 27694 29640 27746 29646
rect 27694 29582 27746 29588
rect 27602 28756 27654 28762
rect 27602 28698 27654 28704
rect 27706 26330 27734 29582
rect 27706 26302 27826 26330
rect 27798 18766 27826 26302
rect 27602 18760 27654 18766
rect 27602 18702 27654 18708
rect 27786 18760 27838 18766
rect 27786 18702 27838 18708
rect 27510 4140 27562 4146
rect 27510 4082 27562 4088
rect 27510 3732 27562 3738
rect 27430 3692 27510 3720
rect 27510 3674 27562 3680
rect 27418 3052 27470 3058
rect 27418 2994 27470 3000
rect 27430 800 27458 2994
rect 27614 800 27642 18702
rect 27890 3058 27918 30874
rect 27970 17876 28022 17882
rect 27970 17818 28022 17824
rect 27982 17610 28010 17818
rect 27970 17604 28022 17610
rect 27970 17546 28022 17552
rect 28258 8634 28286 55218
rect 29730 53666 29758 56238
rect 29810 55956 29862 55962
rect 29810 55898 29862 55904
rect 29638 53638 29758 53666
rect 28890 50856 28942 50862
rect 28890 50798 28942 50804
rect 28338 41064 28390 41070
rect 28338 41006 28390 41012
rect 28246 8628 28298 8634
rect 28246 8570 28298 8576
rect 28154 4004 28206 4010
rect 28154 3946 28206 3952
rect 27878 3052 27930 3058
rect 27878 2994 27930 3000
rect 27786 2644 27838 2650
rect 27786 2586 27838 2592
rect 27798 800 27826 2586
rect 28166 800 28194 3946
rect 28350 3398 28378 41006
rect 28798 40112 28850 40118
rect 28798 40054 28850 40060
rect 28430 31136 28482 31142
rect 28430 31078 28482 31084
rect 28442 27674 28470 31078
rect 28706 30864 28758 30870
rect 28706 30806 28758 30812
rect 28430 27668 28482 27674
rect 28430 27610 28482 27616
rect 28430 24336 28482 24342
rect 28430 24278 28482 24284
rect 28338 3392 28390 3398
rect 28338 3334 28390 3340
rect 28338 3052 28390 3058
rect 28338 2994 28390 3000
rect 28350 800 28378 2994
rect 28442 2922 28470 24278
rect 28522 4140 28574 4146
rect 28522 4082 28574 4088
rect 28430 2916 28482 2922
rect 28430 2858 28482 2864
rect 28534 800 28562 4082
rect 28718 800 28746 30806
rect 28810 3890 28838 40054
rect 28902 4078 28930 50798
rect 29350 48340 29402 48346
rect 29350 48282 29402 48288
rect 29362 38729 29390 48282
rect 29442 45416 29494 45422
rect 29442 45358 29494 45364
rect 29348 38720 29404 38729
rect 29348 38655 29404 38664
rect 29256 38584 29312 38593
rect 29256 38519 29312 38528
rect 28982 38208 29034 38214
rect 28982 38150 29034 38156
rect 28994 7546 29022 38150
rect 29166 27668 29218 27674
rect 29166 27610 29218 27616
rect 29178 14498 29206 27610
rect 29270 24154 29298 38519
rect 29270 24126 29390 24154
rect 29178 14470 29298 14498
rect 29270 9602 29298 14470
rect 29178 9574 29298 9602
rect 28982 7540 29034 7546
rect 28982 7482 29034 7488
rect 28890 4072 28942 4078
rect 28890 4014 28942 4020
rect 28810 3862 28930 3890
rect 28902 800 28930 3862
rect 28994 3738 29114 3754
rect 28982 3732 29114 3738
rect 29034 3726 29114 3732
rect 28982 3674 29034 3680
rect 29086 1902 29114 3726
rect 29074 1896 29126 1902
rect 29074 1838 29126 1844
rect 29178 950 29206 9574
rect 29362 9178 29390 24126
rect 29350 9172 29402 9178
rect 29350 9114 29402 9120
rect 29454 2990 29482 45358
rect 29534 30184 29586 30190
rect 29534 30126 29586 30132
rect 29546 3058 29574 30126
rect 29638 26790 29666 53638
rect 29626 26784 29678 26790
rect 29626 26726 29678 26732
rect 29626 14952 29678 14958
rect 29626 14894 29678 14900
rect 29638 4146 29666 14894
rect 29822 10810 29850 55898
rect 30190 48346 30218 59200
rect 30270 55344 30322 55350
rect 30270 55286 30322 55292
rect 30178 48340 30230 48346
rect 30178 48282 30230 48288
rect 29902 44328 29954 44334
rect 29902 44270 29954 44276
rect 29914 37330 29942 44270
rect 30282 43722 30310 55286
rect 30650 53786 30678 59200
rect 31202 56438 31230 59200
rect 31926 56500 31978 56506
rect 31926 56442 31978 56448
rect 31190 56432 31242 56438
rect 31190 56374 31242 56380
rect 31478 56358 31690 56386
rect 31098 55616 31150 55622
rect 31190 55616 31242 55622
rect 31098 55558 31150 55564
rect 31188 55584 31190 55593
rect 31242 55584 31244 55593
rect 30914 55412 30966 55418
rect 30914 55354 30966 55360
rect 30926 55146 30954 55354
rect 31110 55350 31138 55558
rect 31188 55519 31244 55528
rect 31478 55418 31506 56358
rect 31662 56234 31690 56358
rect 31558 56228 31610 56234
rect 31558 56170 31610 56176
rect 31650 56228 31702 56234
rect 31650 56170 31702 56176
rect 31570 55729 31598 56170
rect 31648 56128 31704 56137
rect 31648 56063 31704 56072
rect 31832 56128 31888 56137
rect 31832 56063 31888 56072
rect 31662 55962 31690 56063
rect 31650 55956 31702 55962
rect 31650 55898 31702 55904
rect 31742 55956 31794 55962
rect 31742 55898 31794 55904
rect 31754 55729 31782 55898
rect 31556 55720 31612 55729
rect 31556 55655 31612 55664
rect 31740 55720 31796 55729
rect 31740 55655 31796 55664
rect 31846 55418 31874 56063
rect 31938 55690 31966 56442
rect 31926 55684 31978 55690
rect 31926 55626 31978 55632
rect 32018 55684 32070 55690
rect 32018 55626 32070 55632
rect 31466 55412 31518 55418
rect 31466 55354 31518 55360
rect 31834 55412 31886 55418
rect 31834 55354 31886 55360
rect 32030 55350 32058 55626
rect 31098 55344 31150 55350
rect 31098 55286 31150 55292
rect 32018 55344 32070 55350
rect 32018 55286 32070 55292
rect 32214 55282 32242 59200
rect 32476 56264 32532 56273
rect 32476 56199 32532 56208
rect 32202 55276 32254 55282
rect 32202 55218 32254 55224
rect 31006 55208 31058 55214
rect 31006 55150 31058 55156
rect 32386 55208 32438 55214
rect 32386 55150 32438 55156
rect 30914 55140 30966 55146
rect 30914 55082 30966 55088
rect 30638 53780 30690 53786
rect 30638 53722 30690 53728
rect 30270 43716 30322 43722
rect 30270 43658 30322 43664
rect 29902 37324 29954 37330
rect 29902 37266 29954 37272
rect 29994 37324 30046 37330
rect 29994 37266 30046 37272
rect 30006 14498 30034 37266
rect 30006 14470 30126 14498
rect 29810 10804 29862 10810
rect 29810 10746 29862 10752
rect 29994 7540 30046 7546
rect 29994 7482 30046 7488
rect 29626 4140 29678 4146
rect 29626 4082 29678 4088
rect 29626 3120 29678 3126
rect 29626 3062 29678 3068
rect 29534 3052 29586 3058
rect 29534 2994 29586 3000
rect 29350 2984 29402 2990
rect 29350 2926 29402 2932
rect 29442 2984 29494 2990
rect 29442 2926 29494 2932
rect 29362 1426 29390 2926
rect 29350 1420 29402 1426
rect 29350 1362 29402 1368
rect 29166 944 29218 950
rect 29166 886 29218 892
rect 29258 944 29310 950
rect 29258 886 29310 892
rect 29270 800 29298 886
rect 29638 800 29666 3062
rect 30006 800 30034 7482
rect 30098 4690 30126 14470
rect 31018 9450 31046 55150
rect 31650 26308 31702 26314
rect 31650 26250 31702 26256
rect 31558 25152 31610 25158
rect 31558 25094 31610 25100
rect 31570 14498 31598 25094
rect 31294 14470 31598 14498
rect 31006 9444 31058 9450
rect 31006 9386 31058 9392
rect 31006 7540 31058 7546
rect 31006 7482 31058 7488
rect 30086 4684 30138 4690
rect 30086 4626 30138 4632
rect 30178 4072 30230 4078
rect 30178 4014 30230 4020
rect 30190 2038 30218 4014
rect 30822 2848 30874 2854
rect 30822 2790 30874 2796
rect 30834 2650 30862 2790
rect 30822 2644 30874 2650
rect 30822 2586 30874 2592
rect 30638 2100 30690 2106
rect 30638 2042 30690 2048
rect 30178 2032 30230 2038
rect 30178 1974 30230 1980
rect 30270 1420 30322 1426
rect 30270 1362 30322 1368
rect 30282 800 30310 1362
rect 30650 800 30678 2042
rect 31018 800 31046 7482
rect 31098 3392 31150 3398
rect 31098 3334 31150 3340
rect 31110 2922 31138 3334
rect 31098 2916 31150 2922
rect 31098 2858 31150 2864
rect 31294 2106 31322 14470
rect 31662 7562 31690 26250
rect 32110 24200 32162 24206
rect 32110 24142 32162 24148
rect 31386 7534 31690 7562
rect 31282 2100 31334 2106
rect 31282 2042 31334 2048
rect 31386 800 31414 7534
rect 31650 4548 31702 4554
rect 31650 4490 31702 4496
rect 31662 4146 31690 4490
rect 31834 4480 31886 4486
rect 31834 4422 31886 4428
rect 31650 4140 31702 4146
rect 31650 4082 31702 4088
rect 31846 3942 31874 4422
rect 31742 3936 31794 3942
rect 31740 3904 31742 3913
rect 31834 3936 31886 3942
rect 31794 3904 31796 3913
rect 31834 3878 31886 3884
rect 31740 3839 31796 3848
rect 31742 3732 31794 3738
rect 31742 3674 31794 3680
rect 31650 3528 31702 3534
rect 31650 3470 31702 3476
rect 31662 3398 31690 3470
rect 31650 3392 31702 3398
rect 31650 3334 31702 3340
rect 31754 800 31782 3674
rect 31834 3664 31886 3670
rect 31834 3606 31886 3612
rect 31846 3369 31874 3606
rect 31832 3360 31888 3369
rect 31832 3295 31888 3304
rect 32122 800 32150 24142
rect 32398 13938 32426 55150
rect 32490 32774 32518 56199
rect 32766 55350 32794 59200
rect 32938 56296 32990 56302
rect 32938 56238 32990 56244
rect 33030 56296 33082 56302
rect 33030 56238 33082 56244
rect 32950 55978 32978 56238
rect 33042 56166 33070 56238
rect 33214 56228 33266 56234
rect 33214 56170 33266 56176
rect 33030 56160 33082 56166
rect 33030 56102 33082 56108
rect 32950 55950 33162 55978
rect 33226 55962 33254 56170
rect 32938 55412 32990 55418
rect 32938 55354 32990 55360
rect 32754 55344 32806 55350
rect 32754 55286 32806 55292
rect 32950 55146 32978 55354
rect 33030 55276 33082 55282
rect 33030 55218 33082 55224
rect 32938 55140 32990 55146
rect 32938 55082 32990 55088
rect 32478 32768 32530 32774
rect 32478 32710 32530 32716
rect 32938 26376 32990 26382
rect 32938 26318 32990 26324
rect 32478 23588 32530 23594
rect 32478 23530 32530 23536
rect 32386 13932 32438 13938
rect 32386 13874 32438 13880
rect 32294 9920 32346 9926
rect 32294 9862 32346 9868
rect 32306 9722 32334 9862
rect 32294 9716 32346 9722
rect 32294 9658 32346 9664
rect 32490 3777 32518 23530
rect 32846 4004 32898 4010
rect 32846 3946 32898 3952
rect 32476 3768 32532 3777
rect 32476 3703 32532 3712
rect 32478 2644 32530 2650
rect 32478 2586 32530 2592
rect 32490 800 32518 2586
rect 32858 800 32886 3946
rect 32950 3738 32978 26318
rect 33042 22642 33070 55218
rect 33134 55196 33162 55950
rect 33214 55956 33266 55962
rect 33214 55898 33266 55904
rect 33214 55208 33266 55214
rect 33134 55168 33214 55196
rect 33214 55150 33266 55156
rect 33030 22636 33082 22642
rect 33030 22578 33082 22584
rect 33214 18148 33266 18154
rect 33214 18090 33266 18096
rect 33122 17332 33174 17338
rect 33226 17320 33254 18090
rect 33174 17292 33254 17320
rect 33122 17274 33174 17280
rect 33318 11014 33346 59200
rect 33764 56400 33820 56409
rect 33764 56335 33820 56344
rect 33778 22166 33806 56335
rect 33870 55758 33898 59200
rect 33858 55752 33910 55758
rect 33858 55694 33910 55700
rect 33950 55752 34002 55758
rect 33950 55694 34002 55700
rect 33962 55282 33990 55694
rect 33950 55276 34002 55282
rect 33950 55218 34002 55224
rect 33858 55072 33910 55078
rect 33858 55014 33910 55020
rect 33870 43110 33898 55014
rect 34042 48680 34094 48686
rect 34042 48622 34094 48628
rect 33858 43104 33910 43110
rect 33858 43046 33910 43052
rect 33766 22160 33818 22166
rect 33766 22102 33818 22108
rect 33306 11008 33358 11014
rect 33306 10950 33358 10956
rect 33950 4072 34002 4078
rect 33950 4014 34002 4020
rect 33214 3936 33266 3942
rect 33028 3904 33084 3913
rect 33214 3878 33266 3884
rect 33028 3839 33084 3848
rect 33042 3738 33070 3839
rect 32938 3732 32990 3738
rect 32938 3674 32990 3680
rect 33030 3732 33082 3738
rect 33030 3674 33082 3680
rect 33226 800 33254 3878
rect 33672 3360 33728 3369
rect 33672 3295 33728 3304
rect 33686 2922 33714 3295
rect 33582 2916 33634 2922
rect 33582 2858 33634 2864
rect 33674 2916 33726 2922
rect 33674 2858 33726 2864
rect 33594 800 33622 2858
rect 33962 800 33990 4014
rect 34054 3777 34082 48622
rect 34330 36786 34358 59200
rect 34882 57866 34910 59200
rect 34686 57860 34738 57866
rect 34686 57802 34738 57808
rect 34870 57860 34922 57866
rect 34870 57802 34922 57808
rect 34698 48346 34726 57802
rect 34922 57692 35218 57712
rect 34978 57690 35002 57692
rect 35058 57690 35082 57692
rect 35138 57690 35162 57692
rect 35000 57638 35002 57690
rect 35064 57638 35076 57690
rect 35138 57638 35140 57690
rect 34978 57636 35002 57638
rect 35058 57636 35082 57638
rect 35138 57636 35162 57638
rect 34922 57616 35218 57636
rect 34922 56604 35218 56624
rect 34978 56602 35002 56604
rect 35058 56602 35082 56604
rect 35138 56602 35162 56604
rect 35000 56550 35002 56602
rect 35064 56550 35076 56602
rect 35138 56550 35140 56602
rect 34978 56548 35002 56550
rect 35058 56548 35082 56550
rect 35138 56548 35162 56550
rect 34922 56528 35218 56548
rect 35434 56114 35462 59200
rect 35894 56370 35922 59200
rect 35974 56500 36026 56506
rect 35974 56442 36026 56448
rect 36066 56500 36118 56506
rect 36066 56442 36118 56448
rect 35986 56370 36014 56442
rect 35882 56364 35934 56370
rect 35882 56306 35934 56312
rect 35974 56364 36026 56370
rect 35974 56306 36026 56312
rect 36078 56302 36106 56442
rect 36526 56364 36578 56370
rect 36526 56306 36578 56312
rect 36066 56296 36118 56302
rect 36066 56238 36118 56244
rect 35342 56086 35462 56114
rect 35342 55690 35370 56086
rect 35422 55956 35474 55962
rect 35422 55898 35474 55904
rect 35330 55684 35382 55690
rect 35330 55626 35382 55632
rect 34922 55516 35218 55536
rect 34978 55514 35002 55516
rect 35058 55514 35082 55516
rect 35138 55514 35162 55516
rect 35000 55462 35002 55514
rect 35064 55462 35076 55514
rect 35138 55462 35140 55514
rect 34978 55460 35002 55462
rect 35058 55460 35082 55462
rect 35138 55460 35162 55462
rect 34922 55440 35218 55460
rect 35330 55276 35382 55282
rect 35330 55218 35382 55224
rect 34922 54428 35218 54448
rect 34978 54426 35002 54428
rect 35058 54426 35082 54428
rect 35138 54426 35162 54428
rect 35000 54374 35002 54426
rect 35064 54374 35076 54426
rect 35138 54374 35140 54426
rect 34978 54372 35002 54374
rect 35058 54372 35082 54374
rect 35138 54372 35162 54374
rect 34922 54352 35218 54372
rect 34922 53340 35218 53360
rect 34978 53338 35002 53340
rect 35058 53338 35082 53340
rect 35138 53338 35162 53340
rect 35000 53286 35002 53338
rect 35064 53286 35076 53338
rect 35138 53286 35140 53338
rect 34978 53284 35002 53286
rect 35058 53284 35082 53286
rect 35138 53284 35162 53286
rect 34922 53264 35218 53284
rect 34922 52252 35218 52272
rect 34978 52250 35002 52252
rect 35058 52250 35082 52252
rect 35138 52250 35162 52252
rect 35000 52198 35002 52250
rect 35064 52198 35076 52250
rect 35138 52198 35140 52250
rect 34978 52196 35002 52198
rect 35058 52196 35082 52198
rect 35138 52196 35162 52198
rect 34922 52176 35218 52196
rect 34922 51164 35218 51184
rect 34978 51162 35002 51164
rect 35058 51162 35082 51164
rect 35138 51162 35162 51164
rect 35000 51110 35002 51162
rect 35064 51110 35076 51162
rect 35138 51110 35140 51162
rect 34978 51108 35002 51110
rect 35058 51108 35082 51110
rect 35138 51108 35162 51110
rect 34922 51088 35218 51108
rect 34922 50076 35218 50096
rect 34978 50074 35002 50076
rect 35058 50074 35082 50076
rect 35138 50074 35162 50076
rect 35000 50022 35002 50074
rect 35064 50022 35076 50074
rect 35138 50022 35140 50074
rect 34978 50020 35002 50022
rect 35058 50020 35082 50022
rect 35138 50020 35162 50022
rect 34922 50000 35218 50020
rect 34922 48988 35218 49008
rect 34978 48986 35002 48988
rect 35058 48986 35082 48988
rect 35138 48986 35162 48988
rect 35000 48934 35002 48986
rect 35064 48934 35076 48986
rect 35138 48934 35140 48986
rect 34978 48932 35002 48934
rect 35058 48932 35082 48934
rect 35138 48932 35162 48934
rect 34922 48912 35218 48932
rect 34594 48340 34646 48346
rect 34594 48282 34646 48288
rect 34686 48340 34738 48346
rect 34686 48282 34738 48288
rect 34410 48000 34462 48006
rect 34410 47942 34462 47948
rect 34318 36780 34370 36786
rect 34318 36722 34370 36728
rect 34422 4078 34450 47942
rect 34606 43382 34634 48282
rect 34922 47900 35218 47920
rect 34978 47898 35002 47900
rect 35058 47898 35082 47900
rect 35138 47898 35162 47900
rect 35000 47846 35002 47898
rect 35064 47846 35076 47898
rect 35138 47846 35140 47898
rect 34978 47844 35002 47846
rect 35058 47844 35082 47846
rect 35138 47844 35162 47846
rect 34922 47824 35218 47844
rect 34922 46812 35218 46832
rect 34978 46810 35002 46812
rect 35058 46810 35082 46812
rect 35138 46810 35162 46812
rect 35000 46758 35002 46810
rect 35064 46758 35076 46810
rect 35138 46758 35140 46810
rect 34978 46756 35002 46758
rect 35058 46756 35082 46758
rect 35138 46756 35162 46758
rect 34922 46736 35218 46756
rect 34922 45724 35218 45744
rect 34978 45722 35002 45724
rect 35058 45722 35082 45724
rect 35138 45722 35162 45724
rect 35000 45670 35002 45722
rect 35064 45670 35076 45722
rect 35138 45670 35140 45722
rect 34978 45668 35002 45670
rect 35058 45668 35082 45670
rect 35138 45668 35162 45670
rect 34922 45648 35218 45668
rect 34922 44636 35218 44656
rect 34978 44634 35002 44636
rect 35058 44634 35082 44636
rect 35138 44634 35162 44636
rect 35000 44582 35002 44634
rect 35064 44582 35076 44634
rect 35138 44582 35140 44634
rect 34978 44580 35002 44582
rect 35058 44580 35082 44582
rect 35138 44580 35162 44582
rect 34922 44560 35218 44580
rect 34922 43548 35218 43568
rect 34978 43546 35002 43548
rect 35058 43546 35082 43548
rect 35138 43546 35162 43548
rect 35000 43494 35002 43546
rect 35064 43494 35076 43546
rect 35138 43494 35140 43546
rect 34978 43492 35002 43494
rect 35058 43492 35082 43494
rect 35138 43492 35162 43494
rect 34922 43472 35218 43492
rect 34594 43376 34646 43382
rect 34594 43318 34646 43324
rect 34778 43376 34830 43382
rect 34778 43318 34830 43324
rect 34790 29034 34818 43318
rect 34922 42460 35218 42480
rect 34978 42458 35002 42460
rect 35058 42458 35082 42460
rect 35138 42458 35162 42460
rect 35000 42406 35002 42458
rect 35064 42406 35076 42458
rect 35138 42406 35140 42458
rect 34978 42404 35002 42406
rect 35058 42404 35082 42406
rect 35138 42404 35162 42406
rect 34922 42384 35218 42404
rect 34922 41372 35218 41392
rect 34978 41370 35002 41372
rect 35058 41370 35082 41372
rect 35138 41370 35162 41372
rect 35000 41318 35002 41370
rect 35064 41318 35076 41370
rect 35138 41318 35140 41370
rect 34978 41316 35002 41318
rect 35058 41316 35082 41318
rect 35138 41316 35162 41318
rect 34922 41296 35218 41316
rect 34922 40284 35218 40304
rect 34978 40282 35002 40284
rect 35058 40282 35082 40284
rect 35138 40282 35162 40284
rect 35000 40230 35002 40282
rect 35064 40230 35076 40282
rect 35138 40230 35140 40282
rect 34978 40228 35002 40230
rect 35058 40228 35082 40230
rect 35138 40228 35162 40230
rect 34922 40208 35218 40228
rect 34922 39196 35218 39216
rect 34978 39194 35002 39196
rect 35058 39194 35082 39196
rect 35138 39194 35162 39196
rect 35000 39142 35002 39194
rect 35064 39142 35076 39194
rect 35138 39142 35140 39194
rect 34978 39140 35002 39142
rect 35058 39140 35082 39142
rect 35138 39140 35162 39142
rect 34922 39120 35218 39140
rect 34922 38108 35218 38128
rect 34978 38106 35002 38108
rect 35058 38106 35082 38108
rect 35138 38106 35162 38108
rect 35000 38054 35002 38106
rect 35064 38054 35076 38106
rect 35138 38054 35140 38106
rect 34978 38052 35002 38054
rect 35058 38052 35082 38054
rect 35138 38052 35162 38054
rect 34922 38032 35218 38052
rect 34922 37020 35218 37040
rect 34978 37018 35002 37020
rect 35058 37018 35082 37020
rect 35138 37018 35162 37020
rect 35000 36966 35002 37018
rect 35064 36966 35076 37018
rect 35138 36966 35140 37018
rect 34978 36964 35002 36966
rect 35058 36964 35082 36966
rect 35138 36964 35162 36966
rect 34922 36944 35218 36964
rect 35238 36712 35290 36718
rect 35238 36654 35290 36660
rect 34922 35932 35218 35952
rect 34978 35930 35002 35932
rect 35058 35930 35082 35932
rect 35138 35930 35162 35932
rect 35000 35878 35002 35930
rect 35064 35878 35076 35930
rect 35138 35878 35140 35930
rect 34978 35876 35002 35878
rect 35058 35876 35082 35878
rect 35138 35876 35162 35878
rect 34922 35856 35218 35876
rect 34922 34844 35218 34864
rect 34978 34842 35002 34844
rect 35058 34842 35082 34844
rect 35138 34842 35162 34844
rect 35000 34790 35002 34842
rect 35064 34790 35076 34842
rect 35138 34790 35140 34842
rect 34978 34788 35002 34790
rect 35058 34788 35082 34790
rect 35138 34788 35162 34790
rect 34922 34768 35218 34788
rect 34922 33756 35218 33776
rect 34978 33754 35002 33756
rect 35058 33754 35082 33756
rect 35138 33754 35162 33756
rect 35000 33702 35002 33754
rect 35064 33702 35076 33754
rect 35138 33702 35140 33754
rect 34978 33700 35002 33702
rect 35058 33700 35082 33702
rect 35138 33700 35162 33702
rect 34922 33680 35218 33700
rect 34922 32668 35218 32688
rect 34978 32666 35002 32668
rect 35058 32666 35082 32668
rect 35138 32666 35162 32668
rect 35000 32614 35002 32666
rect 35064 32614 35076 32666
rect 35138 32614 35140 32666
rect 34978 32612 35002 32614
rect 35058 32612 35082 32614
rect 35138 32612 35162 32614
rect 34922 32592 35218 32612
rect 34922 31580 35218 31600
rect 34978 31578 35002 31580
rect 35058 31578 35082 31580
rect 35138 31578 35162 31580
rect 35000 31526 35002 31578
rect 35064 31526 35076 31578
rect 35138 31526 35140 31578
rect 34978 31524 35002 31526
rect 35058 31524 35082 31526
rect 35138 31524 35162 31526
rect 34922 31504 35218 31524
rect 34922 30492 35218 30512
rect 34978 30490 35002 30492
rect 35058 30490 35082 30492
rect 35138 30490 35162 30492
rect 35000 30438 35002 30490
rect 35064 30438 35076 30490
rect 35138 30438 35140 30490
rect 34978 30436 35002 30438
rect 35058 30436 35082 30438
rect 35138 30436 35162 30438
rect 34922 30416 35218 30436
rect 34922 29404 35218 29424
rect 34978 29402 35002 29404
rect 35058 29402 35082 29404
rect 35138 29402 35162 29404
rect 35000 29350 35002 29402
rect 35064 29350 35076 29402
rect 35138 29350 35140 29402
rect 34978 29348 35002 29350
rect 35058 29348 35082 29350
rect 35138 29348 35162 29350
rect 34922 29328 35218 29348
rect 34686 29028 34738 29034
rect 34686 28970 34738 28976
rect 34778 29028 34830 29034
rect 34778 28970 34830 28976
rect 34698 24154 34726 28970
rect 34778 28416 34830 28422
rect 34778 28358 34830 28364
rect 34790 28218 34818 28358
rect 34922 28316 35218 28336
rect 34978 28314 35002 28316
rect 35058 28314 35082 28316
rect 35138 28314 35162 28316
rect 35000 28262 35002 28314
rect 35064 28262 35076 28314
rect 35138 28262 35140 28314
rect 34978 28260 35002 28262
rect 35058 28260 35082 28262
rect 35138 28260 35162 28262
rect 34922 28240 35218 28260
rect 34778 28212 34830 28218
rect 34778 28154 34830 28160
rect 34922 27228 35218 27248
rect 34978 27226 35002 27228
rect 35058 27226 35082 27228
rect 35138 27226 35162 27228
rect 35000 27174 35002 27226
rect 35064 27174 35076 27226
rect 35138 27174 35140 27226
rect 34978 27172 35002 27174
rect 35058 27172 35082 27174
rect 35138 27172 35162 27174
rect 34922 27152 35218 27172
rect 34922 26140 35218 26160
rect 34978 26138 35002 26140
rect 35058 26138 35082 26140
rect 35138 26138 35162 26140
rect 35000 26086 35002 26138
rect 35064 26086 35076 26138
rect 35138 26086 35140 26138
rect 34978 26084 35002 26086
rect 35058 26084 35082 26086
rect 35138 26084 35162 26086
rect 34922 26064 35218 26084
rect 34922 25052 35218 25072
rect 34978 25050 35002 25052
rect 35058 25050 35082 25052
rect 35138 25050 35162 25052
rect 35000 24998 35002 25050
rect 35064 24998 35076 25050
rect 35138 24998 35140 25050
rect 34978 24996 35002 24998
rect 35058 24996 35082 24998
rect 35138 24996 35162 24998
rect 34922 24976 35218 24996
rect 34606 24126 34726 24154
rect 34606 17218 34634 24126
rect 34922 23964 35218 23984
rect 34978 23962 35002 23964
rect 35058 23962 35082 23964
rect 35138 23962 35162 23964
rect 35000 23910 35002 23962
rect 35064 23910 35076 23962
rect 35138 23910 35140 23962
rect 34978 23908 35002 23910
rect 35058 23908 35082 23910
rect 35138 23908 35162 23910
rect 34922 23888 35218 23908
rect 34922 22876 35218 22896
rect 34978 22874 35002 22876
rect 35058 22874 35082 22876
rect 35138 22874 35162 22876
rect 35000 22822 35002 22874
rect 35064 22822 35076 22874
rect 35138 22822 35140 22874
rect 34978 22820 35002 22822
rect 35058 22820 35082 22822
rect 35138 22820 35162 22822
rect 34922 22800 35218 22820
rect 34922 21788 35218 21808
rect 34978 21786 35002 21788
rect 35058 21786 35082 21788
rect 35138 21786 35162 21788
rect 35000 21734 35002 21786
rect 35064 21734 35076 21786
rect 35138 21734 35140 21786
rect 34978 21732 35002 21734
rect 35058 21732 35082 21734
rect 35138 21732 35162 21734
rect 34922 21712 35218 21732
rect 34922 20700 35218 20720
rect 34978 20698 35002 20700
rect 35058 20698 35082 20700
rect 35138 20698 35162 20700
rect 35000 20646 35002 20698
rect 35064 20646 35076 20698
rect 35138 20646 35140 20698
rect 34978 20644 35002 20646
rect 35058 20644 35082 20646
rect 35138 20644 35162 20646
rect 34922 20624 35218 20644
rect 34922 19612 35218 19632
rect 34978 19610 35002 19612
rect 35058 19610 35082 19612
rect 35138 19610 35162 19612
rect 35000 19558 35002 19610
rect 35064 19558 35076 19610
rect 35138 19558 35140 19610
rect 34978 19556 35002 19558
rect 35058 19556 35082 19558
rect 35138 19556 35162 19558
rect 34922 19536 35218 19556
rect 34922 18524 35218 18544
rect 34978 18522 35002 18524
rect 35058 18522 35082 18524
rect 35138 18522 35162 18524
rect 35000 18470 35002 18522
rect 35064 18470 35076 18522
rect 35138 18470 35140 18522
rect 34978 18468 35002 18470
rect 35058 18468 35082 18470
rect 35138 18468 35162 18470
rect 34922 18448 35218 18468
rect 34922 17436 35218 17456
rect 34978 17434 35002 17436
rect 35058 17434 35082 17436
rect 35138 17434 35162 17436
rect 35000 17382 35002 17434
rect 35064 17382 35076 17434
rect 35138 17382 35140 17434
rect 34978 17380 35002 17382
rect 35058 17380 35082 17382
rect 35138 17380 35162 17382
rect 34922 17360 35218 17380
rect 34514 17190 34634 17218
rect 34514 10266 34542 17190
rect 34922 16348 35218 16368
rect 34978 16346 35002 16348
rect 35058 16346 35082 16348
rect 35138 16346 35162 16348
rect 35000 16294 35002 16346
rect 35064 16294 35076 16346
rect 35138 16294 35140 16346
rect 34978 16292 35002 16294
rect 35058 16292 35082 16294
rect 35138 16292 35162 16294
rect 34922 16272 35218 16292
rect 34594 16040 34646 16046
rect 34594 15982 34646 15988
rect 34778 16040 34830 16046
rect 34778 15982 34830 15988
rect 34502 10260 34554 10266
rect 34502 10202 34554 10208
rect 34606 4078 34634 15982
rect 34686 7472 34738 7478
rect 34686 7414 34738 7420
rect 34410 4072 34462 4078
rect 34410 4014 34462 4020
rect 34594 4072 34646 4078
rect 34594 4014 34646 4020
rect 34040 3768 34096 3777
rect 34040 3703 34096 3712
rect 34594 3392 34646 3398
rect 34594 3334 34646 3340
rect 34500 3224 34556 3233
rect 34500 3159 34556 3168
rect 34514 2961 34542 3159
rect 34500 2952 34556 2961
rect 34606 2922 34634 3334
rect 34500 2887 34556 2896
rect 34594 2916 34646 2922
rect 34594 2858 34646 2864
rect 34318 2848 34370 2854
rect 34318 2790 34370 2796
rect 34330 800 34358 2790
rect 34698 800 34726 7414
rect 34790 1986 34818 15982
rect 34922 15260 35218 15280
rect 34978 15258 35002 15260
rect 35058 15258 35082 15260
rect 35138 15258 35162 15260
rect 35000 15206 35002 15258
rect 35064 15206 35076 15258
rect 35138 15206 35140 15258
rect 34978 15204 35002 15206
rect 35058 15204 35082 15206
rect 35138 15204 35162 15206
rect 34922 15184 35218 15204
rect 34922 14172 35218 14192
rect 34978 14170 35002 14172
rect 35058 14170 35082 14172
rect 35138 14170 35162 14172
rect 35000 14118 35002 14170
rect 35064 14118 35076 14170
rect 35138 14118 35140 14170
rect 34978 14116 35002 14118
rect 35058 14116 35082 14118
rect 35138 14116 35162 14118
rect 34922 14096 35218 14116
rect 34922 13084 35218 13104
rect 34978 13082 35002 13084
rect 35058 13082 35082 13084
rect 35138 13082 35162 13084
rect 35000 13030 35002 13082
rect 35064 13030 35076 13082
rect 35138 13030 35140 13082
rect 34978 13028 35002 13030
rect 35058 13028 35082 13030
rect 35138 13028 35162 13030
rect 34922 13008 35218 13028
rect 34922 11996 35218 12016
rect 34978 11994 35002 11996
rect 35058 11994 35082 11996
rect 35138 11994 35162 11996
rect 35000 11942 35002 11994
rect 35064 11942 35076 11994
rect 35138 11942 35140 11994
rect 34978 11940 35002 11942
rect 35058 11940 35082 11942
rect 35138 11940 35162 11942
rect 34922 11920 35218 11940
rect 34922 10908 35218 10928
rect 34978 10906 35002 10908
rect 35058 10906 35082 10908
rect 35138 10906 35162 10908
rect 35000 10854 35002 10906
rect 35064 10854 35076 10906
rect 35138 10854 35140 10906
rect 34978 10852 35002 10854
rect 35058 10852 35082 10854
rect 35138 10852 35162 10854
rect 34922 10832 35218 10852
rect 34922 9820 35218 9840
rect 34978 9818 35002 9820
rect 35058 9818 35082 9820
rect 35138 9818 35162 9820
rect 35000 9766 35002 9818
rect 35064 9766 35076 9818
rect 35138 9766 35140 9818
rect 34978 9764 35002 9766
rect 35058 9764 35082 9766
rect 35138 9764 35162 9766
rect 34922 9744 35218 9764
rect 34922 8732 35218 8752
rect 34978 8730 35002 8732
rect 35058 8730 35082 8732
rect 35138 8730 35162 8732
rect 35000 8678 35002 8730
rect 35064 8678 35076 8730
rect 35138 8678 35140 8730
rect 34978 8676 35002 8678
rect 35058 8676 35082 8678
rect 35138 8676 35162 8678
rect 34922 8656 35218 8676
rect 34922 7644 35218 7664
rect 34978 7642 35002 7644
rect 35058 7642 35082 7644
rect 35138 7642 35162 7644
rect 35000 7590 35002 7642
rect 35064 7590 35076 7642
rect 35138 7590 35140 7642
rect 34978 7588 35002 7590
rect 35058 7588 35082 7590
rect 35138 7588 35162 7590
rect 34922 7568 35218 7588
rect 34922 6556 35218 6576
rect 34978 6554 35002 6556
rect 35058 6554 35082 6556
rect 35138 6554 35162 6556
rect 35000 6502 35002 6554
rect 35064 6502 35076 6554
rect 35138 6502 35140 6554
rect 34978 6500 35002 6502
rect 35058 6500 35082 6502
rect 35138 6500 35162 6502
rect 34922 6480 35218 6500
rect 34922 5468 35218 5488
rect 34978 5466 35002 5468
rect 35058 5466 35082 5468
rect 35138 5466 35162 5468
rect 35000 5414 35002 5466
rect 35064 5414 35076 5466
rect 35138 5414 35140 5466
rect 34978 5412 35002 5414
rect 35058 5412 35082 5414
rect 35138 5412 35162 5414
rect 34922 5392 35218 5412
rect 34922 4380 35218 4400
rect 34978 4378 35002 4380
rect 35058 4378 35082 4380
rect 35138 4378 35162 4380
rect 35000 4326 35002 4378
rect 35064 4326 35076 4378
rect 35138 4326 35140 4378
rect 34978 4324 35002 4326
rect 35058 4324 35082 4326
rect 35138 4324 35162 4326
rect 34922 4304 35218 4324
rect 35250 3942 35278 36654
rect 35342 15162 35370 55218
rect 35434 48278 35462 55898
rect 35882 55752 35934 55758
rect 35882 55694 35934 55700
rect 35894 52426 35922 55694
rect 35882 52420 35934 52426
rect 35882 52362 35934 52368
rect 35422 48272 35474 48278
rect 35422 48214 35474 48220
rect 35514 48204 35566 48210
rect 35514 48146 35566 48152
rect 35526 21894 35554 48146
rect 35514 21888 35566 21894
rect 35514 21830 35566 21836
rect 36538 16250 36566 56306
rect 36998 55418 37026 59200
rect 37550 55826 37578 59200
rect 37538 55820 37590 55826
rect 37538 55762 37590 55768
rect 37630 55820 37682 55826
rect 37630 55762 37682 55768
rect 37078 55684 37130 55690
rect 37078 55626 37130 55632
rect 37090 55418 37118 55626
rect 36986 55412 37038 55418
rect 36986 55354 37038 55360
rect 37078 55412 37130 55418
rect 37078 55354 37130 55360
rect 37642 55078 37670 55762
rect 38562 55758 38590 59200
rect 38642 55956 38694 55962
rect 38642 55898 38694 55904
rect 38654 55758 38682 55898
rect 38550 55752 38602 55758
rect 38550 55694 38602 55700
rect 38642 55752 38694 55758
rect 38642 55694 38694 55700
rect 38090 55684 38142 55690
rect 38090 55626 38142 55632
rect 37630 55072 37682 55078
rect 37630 55014 37682 55020
rect 38102 48346 38130 55626
rect 38274 55616 38326 55622
rect 38274 55558 38326 55564
rect 37998 48340 38050 48346
rect 37998 48282 38050 48288
rect 38090 48340 38142 48346
rect 38090 48282 38142 48288
rect 36618 44328 36670 44334
rect 36618 44270 36670 44276
rect 36526 16244 36578 16250
rect 36526 16186 36578 16192
rect 35330 15156 35382 15162
rect 35330 15098 35382 15104
rect 36630 3942 36658 44270
rect 37446 43784 37498 43790
rect 37446 43726 37498 43732
rect 36986 39296 37038 39302
rect 36986 39238 37038 39244
rect 35238 3936 35290 3942
rect 35238 3878 35290 3884
rect 36526 3936 36578 3942
rect 36526 3878 36578 3884
rect 36618 3936 36670 3942
rect 36618 3878 36670 3884
rect 36538 3720 36566 3878
rect 36538 3692 36658 3720
rect 36630 3602 36658 3692
rect 36618 3596 36670 3602
rect 36618 3538 36670 3544
rect 36526 3392 36578 3398
rect 36526 3334 36578 3340
rect 34922 3292 35218 3312
rect 34978 3290 35002 3292
rect 35058 3290 35082 3292
rect 35138 3290 35162 3292
rect 35000 3238 35002 3290
rect 35064 3238 35076 3290
rect 35138 3238 35140 3290
rect 34978 3236 35002 3238
rect 35058 3236 35082 3238
rect 35138 3236 35162 3238
rect 34922 3216 35218 3236
rect 36158 3188 36210 3194
rect 36158 3130 36210 3136
rect 35420 2952 35476 2961
rect 35420 2887 35476 2896
rect 34922 2204 35218 2224
rect 34978 2202 35002 2204
rect 35058 2202 35082 2204
rect 35138 2202 35162 2204
rect 35000 2150 35002 2202
rect 35064 2150 35076 2202
rect 35138 2150 35140 2202
rect 34978 2148 35002 2150
rect 35058 2148 35082 2150
rect 35138 2148 35162 2150
rect 34922 2128 35218 2148
rect 34790 1958 35094 1986
rect 35066 800 35094 1958
rect 35434 800 35462 2887
rect 35790 1896 35842 1902
rect 35790 1838 35842 1844
rect 35802 800 35830 1838
rect 36170 800 36198 3130
rect 36538 3058 36566 3334
rect 36526 3052 36578 3058
rect 36526 2994 36578 3000
rect 36526 2032 36578 2038
rect 36526 1974 36578 1980
rect 36538 800 36566 1974
rect 36998 898 37026 39238
rect 37458 37330 37486 43726
rect 37446 37324 37498 37330
rect 37446 37266 37498 37272
rect 37814 28008 37866 28014
rect 37814 27950 37866 27956
rect 37630 25832 37682 25838
rect 37630 25774 37682 25780
rect 37642 25294 37670 25774
rect 37630 25288 37682 25294
rect 37630 25230 37682 25236
rect 37352 16552 37408 16561
rect 37352 16487 37408 16496
rect 37366 11762 37394 16487
rect 37354 11756 37406 11762
rect 37354 11698 37406 11704
rect 37262 4684 37314 4690
rect 37262 4626 37314 4632
rect 36906 870 37026 898
rect 36906 800 36934 870
rect 37274 800 37302 4626
rect 37826 3534 37854 27950
rect 38010 19378 38038 48282
rect 38182 44328 38234 44334
rect 38182 44270 38234 44276
rect 38090 36032 38142 36038
rect 38090 35974 38142 35980
rect 37906 19372 37958 19378
rect 37906 19314 37958 19320
rect 37998 19372 38050 19378
rect 37998 19314 38050 19320
rect 37918 11558 37946 19314
rect 37906 11552 37958 11558
rect 37906 11494 37958 11500
rect 37998 4072 38050 4078
rect 37998 4014 38050 4020
rect 37814 3528 37866 3534
rect 37814 3470 37866 3476
rect 37628 2816 37684 2825
rect 37628 2751 37684 2760
rect 37642 800 37670 2751
rect 38010 800 38038 4014
rect 38102 3126 38130 35974
rect 38090 3120 38142 3126
rect 38090 3062 38142 3068
rect 38194 3058 38222 44270
rect 38286 43466 38314 55558
rect 39114 55162 39142 59200
rect 39470 56772 39522 56778
rect 39470 56714 39522 56720
rect 39482 55350 39510 56714
rect 39470 55344 39522 55350
rect 39470 55286 39522 55292
rect 38654 55134 39142 55162
rect 38286 43438 38498 43466
rect 38470 41290 38498 43438
rect 38378 41262 38498 41290
rect 38378 35834 38406 41262
rect 38550 37120 38602 37126
rect 38550 37062 38602 37068
rect 38366 35828 38418 35834
rect 38366 35770 38418 35776
rect 38274 17536 38326 17542
rect 38274 17478 38326 17484
rect 38286 4554 38314 17478
rect 38274 4548 38326 4554
rect 38274 4490 38326 4496
rect 38562 4078 38590 37062
rect 38654 10674 38682 55134
rect 39574 53106 39602 59200
rect 40126 56438 40154 59200
rect 40114 56432 40166 56438
rect 40206 56432 40258 56438
rect 40114 56374 40166 56380
rect 40204 56400 40206 56409
rect 40258 56400 40260 56409
rect 40204 56335 40260 56344
rect 40678 56302 40706 59200
rect 41402 56500 41454 56506
rect 41402 56442 41454 56448
rect 41494 56500 41546 56506
rect 41494 56442 41546 56448
rect 41310 56432 41362 56438
rect 41124 56400 41180 56409
rect 41310 56374 41362 56380
rect 41124 56335 41126 56344
rect 41178 56335 41180 56344
rect 41126 56306 41178 56312
rect 40666 56296 40718 56302
rect 40666 56238 40718 56244
rect 40758 56296 40810 56302
rect 41322 56273 41350 56374
rect 40758 56238 40810 56244
rect 41308 56264 41364 56273
rect 40770 56114 40798 56238
rect 41414 56250 41442 56442
rect 41506 56409 41534 56442
rect 41492 56400 41548 56409
rect 41492 56335 41548 56344
rect 41414 56234 41626 56250
rect 41414 56228 41638 56234
rect 41414 56222 41586 56228
rect 41308 56199 41364 56208
rect 41586 56170 41638 56176
rect 41690 56166 41718 59200
rect 40586 56086 40798 56114
rect 41402 56160 41454 56166
rect 41678 56160 41730 56166
rect 41454 56108 41534 56114
rect 41402 56102 41534 56108
rect 41678 56102 41730 56108
rect 41414 56086 41534 56102
rect 39654 55956 39706 55962
rect 39654 55898 39706 55904
rect 39010 53100 39062 53106
rect 39010 53042 39062 53048
rect 39562 53100 39614 53106
rect 39562 53042 39614 53048
rect 39022 45558 39050 53042
rect 39666 52986 39694 55898
rect 40586 55826 40614 56086
rect 40574 55820 40626 55826
rect 40574 55762 40626 55768
rect 40666 55820 40718 55826
rect 40666 55762 40718 55768
rect 39298 52958 39694 52986
rect 38826 45552 38878 45558
rect 38826 45494 38878 45500
rect 39010 45552 39062 45558
rect 39010 45494 39062 45500
rect 38838 44169 38866 45494
rect 38824 44160 38880 44169
rect 38824 44095 38880 44104
rect 38826 31272 38878 31278
rect 38826 31214 38878 31220
rect 38734 26240 38786 26246
rect 38734 26182 38786 26188
rect 38746 16697 38774 26182
rect 38732 16688 38788 16697
rect 38732 16623 38788 16632
rect 38642 10668 38694 10674
rect 38642 10610 38694 10616
rect 38550 4072 38602 4078
rect 38550 4014 38602 4020
rect 38642 3596 38694 3602
rect 38642 3538 38694 3544
rect 38734 3596 38786 3602
rect 38734 3538 38786 3544
rect 38366 3188 38418 3194
rect 38366 3130 38418 3136
rect 38182 3052 38234 3058
rect 38182 2994 38234 3000
rect 38378 800 38406 3130
rect 38654 2961 38682 3538
rect 38640 2952 38696 2961
rect 38640 2887 38696 2896
rect 38746 800 38774 3538
rect 38838 1630 38866 31214
rect 39008 26344 39064 26353
rect 39008 26279 39064 26288
rect 39022 26246 39050 26279
rect 39010 26240 39062 26246
rect 39010 26182 39062 26188
rect 39298 17678 39326 52958
rect 39654 52352 39706 52358
rect 39654 52294 39706 52300
rect 39286 17672 39338 17678
rect 39286 17614 39338 17620
rect 39666 4214 39694 52294
rect 39930 30116 39982 30122
rect 39930 30058 39982 30064
rect 39654 4208 39706 4214
rect 39654 4150 39706 4156
rect 39746 4072 39798 4078
rect 39746 4014 39798 4020
rect 39102 3936 39154 3942
rect 39102 3878 39154 3884
rect 39194 3936 39246 3942
rect 39194 3878 39246 3884
rect 38826 1624 38878 1630
rect 38826 1566 38878 1572
rect 39114 800 39142 3878
rect 39206 3738 39234 3878
rect 39194 3732 39246 3738
rect 39194 3674 39246 3680
rect 39758 3058 39786 4014
rect 39942 3602 39970 30058
rect 40678 18154 40706 55762
rect 41506 55622 41534 56086
rect 42242 55690 42270 59200
rect 42230 55684 42282 55690
rect 42230 55626 42282 55632
rect 41402 55616 41454 55622
rect 41402 55558 41454 55564
rect 41494 55616 41546 55622
rect 41494 55558 41546 55564
rect 41308 55448 41364 55457
rect 41414 55434 41442 55558
rect 41414 55418 41718 55434
rect 41414 55412 41730 55418
rect 41414 55406 41678 55412
rect 41308 55383 41310 55392
rect 41362 55383 41364 55392
rect 41310 55354 41362 55360
rect 41678 55354 41730 55360
rect 41310 55276 41362 55282
rect 41494 55276 41546 55282
rect 41362 55236 41494 55264
rect 41310 55218 41362 55224
rect 41494 55218 41546 55224
rect 42794 53122 42822 59200
rect 43254 56234 43282 59200
rect 43242 56228 43294 56234
rect 43242 56170 43294 56176
rect 43806 55418 43834 59200
rect 44910 56778 44938 59200
rect 44898 56772 44950 56778
rect 44898 56714 44950 56720
rect 45370 56234 45398 59200
rect 45922 59158 45950 59200
rect 45726 59152 45778 59158
rect 45726 59094 45778 59100
rect 45910 59152 45962 59158
rect 45910 59094 45962 59100
rect 44162 56228 44214 56234
rect 44162 56170 44214 56176
rect 45358 56228 45410 56234
rect 45358 56170 45410 56176
rect 45450 56228 45502 56234
rect 45450 56170 45502 56176
rect 44174 55894 44202 56170
rect 44898 56160 44950 56166
rect 44898 56102 44950 56108
rect 44162 55888 44214 55894
rect 44162 55830 44214 55836
rect 44714 55888 44766 55894
rect 44714 55830 44766 55836
rect 44622 55684 44674 55690
rect 44622 55626 44674 55632
rect 43794 55412 43846 55418
rect 43794 55354 43846 55360
rect 43886 55412 43938 55418
rect 43886 55354 43938 55360
rect 43610 55344 43662 55350
rect 43610 55286 43662 55292
rect 42794 53094 42914 53122
rect 42886 50946 42914 53094
rect 42886 50918 43006 50946
rect 40758 36644 40810 36650
rect 40758 36586 40810 36592
rect 40666 18148 40718 18154
rect 40666 18090 40718 18096
rect 40666 14000 40718 14006
rect 40666 13942 40718 13948
rect 40298 12096 40350 12102
rect 40298 12038 40350 12044
rect 40310 8294 40338 12038
rect 40678 8566 40706 13942
rect 40666 8560 40718 8566
rect 40666 8502 40718 8508
rect 40298 8288 40350 8294
rect 40298 8230 40350 8236
rect 40206 4820 40258 4826
rect 40206 4762 40258 4768
rect 39930 3596 39982 3602
rect 39930 3538 39982 3544
rect 39930 3460 39982 3466
rect 39930 3402 39982 3408
rect 39746 3052 39798 3058
rect 39746 2994 39798 3000
rect 39470 2984 39522 2990
rect 39470 2926 39522 2932
rect 39482 800 39510 2926
rect 39838 2916 39890 2922
rect 39838 2858 39890 2864
rect 39850 1766 39878 2858
rect 39942 2650 39970 3402
rect 39930 2644 39982 2650
rect 39930 2586 39982 2592
rect 39838 1760 39890 1766
rect 39838 1702 39890 1708
rect 39838 1624 39890 1630
rect 39838 1566 39890 1572
rect 39850 800 39878 1566
rect 40218 800 40246 4762
rect 40770 3942 40798 36586
rect 42046 33856 42098 33862
rect 42046 33798 42098 33804
rect 41126 9716 41178 9722
rect 41126 9658 41178 9664
rect 41138 4826 41166 9658
rect 41402 8560 41454 8566
rect 41402 8502 41454 8508
rect 41126 4820 41178 4826
rect 41126 4762 41178 4768
rect 41034 4480 41086 4486
rect 41034 4422 41086 4428
rect 40574 3936 40626 3942
rect 40574 3878 40626 3884
rect 40758 3936 40810 3942
rect 40758 3878 40810 3884
rect 40390 3664 40442 3670
rect 40390 3606 40442 3612
rect 40402 2582 40430 3606
rect 40390 2576 40442 2582
rect 40390 2518 40442 2524
rect 40586 800 40614 3878
rect 41046 3194 41074 4422
rect 41034 3188 41086 3194
rect 41034 3130 41086 3136
rect 41310 3188 41362 3194
rect 41310 3130 41362 3136
rect 41322 3074 41350 3130
rect 41230 3058 41350 3074
rect 41414 3058 41442 8502
rect 42058 3670 42086 33798
rect 42978 31770 43006 50918
rect 42886 31742 43006 31770
rect 42138 21480 42190 21486
rect 42138 21422 42190 21428
rect 42046 3664 42098 3670
rect 42046 3606 42098 3612
rect 42044 3088 42100 3097
rect 41218 3052 41350 3058
rect 41270 3046 41350 3052
rect 41402 3052 41454 3058
rect 41218 2994 41270 3000
rect 42044 3023 42100 3032
rect 41402 2994 41454 3000
rect 41124 2952 41180 2961
rect 40770 2910 40982 2938
rect 40770 2854 40798 2910
rect 40758 2848 40810 2854
rect 40758 2790 40810 2796
rect 40850 2848 40902 2854
rect 40850 2790 40902 2796
rect 40862 2650 40890 2790
rect 40850 2644 40902 2650
rect 40850 2586 40902 2592
rect 40954 800 40982 2910
rect 41180 2922 41350 2938
rect 41180 2916 41362 2922
rect 41180 2910 41310 2916
rect 41124 2887 41180 2896
rect 41310 2858 41362 2864
rect 41678 2916 41730 2922
rect 41678 2858 41730 2864
rect 41310 1760 41362 1766
rect 41310 1702 41362 1708
rect 41322 800 41350 1702
rect 41690 800 41718 2858
rect 42058 800 42086 3023
rect 42150 2922 42178 21422
rect 42886 12782 42914 31742
rect 43622 24274 43650 55286
rect 43898 55146 43926 55354
rect 43886 55140 43938 55146
rect 43886 55082 43938 55088
rect 43610 24268 43662 24274
rect 43610 24210 43662 24216
rect 44162 18148 44214 18154
rect 44162 18090 44214 18096
rect 42874 12776 42926 12782
rect 42874 12718 42926 12724
rect 44070 12096 44122 12102
rect 44070 12038 44122 12044
rect 43150 4276 43202 4282
rect 43150 4218 43202 4224
rect 42782 2984 42834 2990
rect 42782 2926 42834 2932
rect 42138 2916 42190 2922
rect 42138 2858 42190 2864
rect 42414 2576 42466 2582
rect 42414 2518 42466 2524
rect 42426 800 42454 2518
rect 42794 800 42822 2926
rect 43162 800 43190 4218
rect 43516 4040 43572 4049
rect 43516 3975 43572 3984
rect 43530 800 43558 3975
rect 44082 898 44110 12038
rect 44174 9722 44202 18090
rect 44634 14482 44662 55626
rect 44622 14476 44674 14482
rect 44622 14418 44674 14424
rect 44726 12986 44754 55830
rect 44910 43994 44938 56102
rect 45462 55457 45490 56170
rect 45448 55448 45504 55457
rect 45448 55383 45504 55392
rect 45738 53825 45766 59094
rect 46474 55418 46502 59200
rect 47026 55622 47054 59200
rect 47014 55616 47066 55622
rect 47014 55558 47066 55564
rect 46462 55412 46514 55418
rect 46462 55354 46514 55360
rect 48038 55162 48066 59200
rect 48590 56234 48618 59200
rect 48578 56228 48630 56234
rect 48578 56170 48630 56176
rect 49050 55162 49078 59200
rect 49602 55298 49630 59200
rect 50154 55350 50182 59200
rect 50282 57148 50578 57168
rect 50338 57146 50362 57148
rect 50418 57146 50442 57148
rect 50498 57146 50522 57148
rect 50360 57094 50362 57146
rect 50424 57094 50436 57146
rect 50498 57094 50500 57146
rect 50338 57092 50362 57094
rect 50418 57092 50442 57094
rect 50498 57092 50522 57094
rect 50282 57072 50578 57092
rect 51166 56438 51194 59200
rect 51244 58032 51300 58041
rect 51244 57967 51300 57976
rect 51154 56432 51206 56438
rect 51154 56374 51206 56380
rect 50282 56060 50578 56080
rect 50338 56058 50362 56060
rect 50418 56058 50442 56060
rect 50498 56058 50522 56060
rect 50360 56006 50362 56058
rect 50424 56006 50436 56058
rect 50498 56006 50500 56058
rect 50338 56004 50362 56006
rect 50418 56004 50442 56006
rect 50498 56004 50522 56006
rect 50282 55984 50578 56004
rect 50142 55344 50194 55350
rect 49602 55270 49906 55298
rect 50142 55286 50194 55292
rect 48038 55134 48250 55162
rect 45540 53816 45596 53825
rect 45540 53751 45596 53760
rect 45724 53816 45780 53825
rect 45724 53751 45780 53760
rect 45554 44198 45582 53751
rect 45542 44192 45594 44198
rect 45542 44134 45594 44140
rect 45726 44192 45778 44198
rect 45726 44134 45778 44140
rect 44898 43988 44950 43994
rect 44898 43930 44950 43936
rect 44990 34536 45042 34542
rect 45738 34513 45766 44134
rect 46278 37324 46330 37330
rect 46278 37266 46330 37272
rect 44990 34478 45042 34484
rect 45540 34504 45596 34513
rect 44806 25288 44858 25294
rect 44806 25230 44858 25236
rect 44714 12980 44766 12986
rect 44714 12922 44766 12928
rect 44162 9716 44214 9722
rect 44162 9658 44214 9664
rect 44620 3768 44676 3777
rect 44620 3703 44676 3712
rect 44254 2848 44306 2854
rect 44254 2790 44306 2796
rect 43898 870 44110 898
rect 43898 800 43926 870
rect 44266 800 44294 2790
rect 44634 800 44662 3703
rect 44818 2922 44846 25230
rect 44806 2916 44858 2922
rect 44806 2858 44858 2864
rect 45002 800 45030 34478
rect 45540 34439 45596 34448
rect 45724 34504 45780 34513
rect 45724 34439 45780 34448
rect 45554 24886 45582 34439
rect 45542 24880 45594 24886
rect 45356 24848 45412 24857
rect 45726 24880 45778 24886
rect 45542 24822 45594 24828
rect 45724 24848 45726 24857
rect 45778 24848 45780 24857
rect 45356 24783 45412 24792
rect 45724 24783 45780 24792
rect 45370 15366 45398 24783
rect 46290 18714 46318 37266
rect 48118 30184 48170 30190
rect 48118 30126 48170 30132
rect 48130 29714 48158 30126
rect 48118 29708 48170 29714
rect 48118 29650 48170 29656
rect 47934 21888 47986 21894
rect 47934 21830 47986 21836
rect 46290 18686 46410 18714
rect 45358 15360 45410 15366
rect 45358 15302 45410 15308
rect 45542 15360 45594 15366
rect 45542 15302 45594 15308
rect 45174 14272 45226 14278
rect 45174 14214 45226 14220
rect 45186 898 45214 14214
rect 45554 13870 45582 15302
rect 45542 13864 45594 13870
rect 45542 13806 45594 13812
rect 46278 7744 46330 7750
rect 46278 7686 46330 7692
rect 46290 7546 46318 7686
rect 46278 7540 46330 7546
rect 46278 7482 46330 7488
rect 45726 3460 45778 3466
rect 45726 3402 45778 3408
rect 45266 3188 45318 3194
rect 45266 3130 45318 3136
rect 45278 2990 45306 3130
rect 45266 2984 45318 2990
rect 45266 2926 45318 2932
rect 45186 870 45398 898
rect 45370 800 45398 870
rect 45738 800 45766 3402
rect 46094 3392 46146 3398
rect 46094 3334 46146 3340
rect 46106 800 46134 3334
rect 46382 898 46410 18686
rect 47474 18624 47526 18630
rect 47474 18566 47526 18572
rect 46830 14952 46882 14958
rect 46830 14894 46882 14900
rect 46738 4140 46790 4146
rect 46738 4082 46790 4088
rect 46750 3346 46778 4082
rect 46842 3466 46870 14894
rect 47290 8288 47342 8294
rect 47290 8230 47342 8236
rect 47014 4548 47066 4554
rect 47014 4490 47066 4496
rect 46922 3664 46974 3670
rect 46922 3606 46974 3612
rect 46830 3460 46882 3466
rect 46830 3402 46882 3408
rect 46750 3318 46870 3346
rect 46382 870 46502 898
rect 46474 800 46502 870
rect 46842 800 46870 3318
rect 46934 3194 46962 3606
rect 47026 3466 47054 4490
rect 47196 3632 47252 3641
rect 47196 3567 47252 3576
rect 47014 3460 47066 3466
rect 47014 3402 47066 3408
rect 46922 3188 46974 3194
rect 46922 3130 46974 3136
rect 47210 800 47238 3567
rect 47302 3534 47330 8230
rect 47486 3670 47514 18566
rect 47474 3664 47526 3670
rect 47474 3606 47526 3612
rect 47946 3602 47974 21830
rect 48118 20596 48170 20602
rect 48118 20538 48170 20544
rect 48130 20398 48158 20538
rect 48118 20392 48170 20398
rect 48118 20334 48170 20340
rect 48222 15366 48250 55134
rect 48498 55134 49078 55162
rect 48302 43988 48354 43994
rect 48302 43930 48354 43936
rect 48314 43858 48342 43930
rect 48302 43852 48354 43858
rect 48302 43794 48354 43800
rect 48498 41018 48526 55134
rect 48946 54324 48998 54330
rect 48946 54266 48998 54272
rect 48406 40990 48526 41018
rect 48406 38570 48434 40990
rect 48406 38542 48526 38570
rect 48498 33862 48526 38542
rect 48486 33856 48538 33862
rect 48486 33798 48538 33804
rect 48670 33856 48722 33862
rect 48670 33798 48722 33804
rect 48486 30184 48538 30190
rect 48486 30126 48538 30132
rect 48498 29782 48526 30126
rect 48486 29776 48538 29782
rect 48486 29718 48538 29724
rect 48682 29034 48710 33798
rect 48302 29028 48354 29034
rect 48302 28970 48354 28976
rect 48670 29028 48722 29034
rect 48670 28970 48722 28976
rect 48314 19281 48342 28970
rect 48300 19272 48356 19281
rect 48300 19207 48356 19216
rect 48392 19136 48448 19145
rect 48392 19071 48448 19080
rect 48210 15360 48262 15366
rect 48210 15302 48262 15308
rect 48406 15026 48434 19071
rect 48762 17536 48814 17542
rect 48762 17478 48814 17484
rect 48394 15020 48446 15026
rect 48394 14962 48446 14968
rect 48774 12374 48802 17478
rect 48762 12368 48814 12374
rect 48762 12310 48814 12316
rect 48394 8832 48446 8838
rect 48394 8774 48446 8780
rect 48406 8634 48434 8774
rect 48394 8628 48446 8634
rect 48394 8570 48446 8576
rect 48958 3942 48986 54266
rect 49590 39296 49642 39302
rect 49590 39238 49642 39244
rect 49038 19848 49090 19854
rect 49038 19790 49090 19796
rect 48946 3936 48998 3942
rect 48946 3878 48998 3884
rect 49050 3738 49078 19790
rect 49222 12368 49274 12374
rect 49222 12310 49274 12316
rect 49234 9625 49262 12310
rect 49220 9616 49276 9625
rect 49220 9551 49276 9560
rect 48670 3732 48722 3738
rect 48670 3674 48722 3680
rect 49038 3732 49090 3738
rect 49038 3674 49090 3680
rect 47934 3596 47986 3602
rect 47934 3538 47986 3544
rect 47290 3528 47342 3534
rect 47290 3470 47342 3476
rect 48302 3528 48354 3534
rect 48354 3488 48434 3516
rect 48302 3470 48354 3476
rect 48406 3482 48434 3488
rect 48406 3454 48526 3482
rect 47566 3392 47618 3398
rect 48392 3360 48448 3369
rect 47566 3334 47618 3340
rect 47578 800 47606 3334
rect 48314 3318 48392 3346
rect 47934 3120 47986 3126
rect 47934 3062 47986 3068
rect 47946 800 47974 3062
rect 48314 800 48342 3318
rect 48392 3295 48448 3304
rect 48498 2582 48526 3454
rect 48486 2576 48538 2582
rect 48486 2518 48538 2524
rect 48682 800 48710 3674
rect 49038 2984 49090 2990
rect 49038 2926 49090 2932
rect 49050 800 49078 2926
rect 49602 898 49630 39238
rect 49878 13802 49906 55270
rect 50282 54972 50578 54992
rect 50338 54970 50362 54972
rect 50418 54970 50442 54972
rect 50498 54970 50522 54972
rect 50360 54918 50362 54970
rect 50424 54918 50436 54970
rect 50498 54918 50500 54970
rect 50338 54916 50362 54918
rect 50418 54916 50442 54918
rect 50498 54916 50522 54918
rect 50282 54896 50578 54916
rect 50282 53884 50578 53904
rect 50338 53882 50362 53884
rect 50418 53882 50442 53884
rect 50498 53882 50522 53884
rect 50360 53830 50362 53882
rect 50424 53830 50436 53882
rect 50498 53830 50500 53882
rect 50338 53828 50362 53830
rect 50418 53828 50442 53830
rect 50498 53828 50522 53830
rect 50282 53808 50578 53828
rect 51258 53122 51286 57967
rect 51718 55282 51746 59200
rect 52270 58041 52298 59200
rect 52256 58032 52312 58041
rect 52256 57967 52312 57976
rect 52730 56370 52758 59200
rect 52718 56364 52770 56370
rect 52718 56306 52770 56312
rect 53282 55758 53310 59200
rect 53270 55752 53322 55758
rect 53270 55694 53322 55700
rect 54386 55690 54414 59200
rect 54846 56506 54874 59200
rect 55398 59106 55426 59200
rect 55214 59078 55426 59106
rect 54834 56500 54886 56506
rect 54834 56442 54886 56448
rect 54374 55684 54426 55690
rect 54374 55626 54426 55632
rect 52442 55616 52494 55622
rect 52442 55558 52494 55564
rect 51706 55276 51758 55282
rect 51706 55218 51758 55224
rect 51166 53094 51286 53122
rect 50282 52796 50578 52816
rect 50338 52794 50362 52796
rect 50418 52794 50442 52796
rect 50498 52794 50522 52796
rect 50360 52742 50362 52794
rect 50424 52742 50436 52794
rect 50498 52742 50500 52794
rect 50338 52740 50362 52742
rect 50418 52740 50442 52742
rect 50498 52740 50522 52742
rect 50282 52720 50578 52740
rect 50282 51708 50578 51728
rect 50338 51706 50362 51708
rect 50418 51706 50442 51708
rect 50498 51706 50522 51708
rect 50360 51654 50362 51706
rect 50424 51654 50436 51706
rect 50498 51654 50500 51706
rect 50338 51652 50362 51654
rect 50418 51652 50442 51654
rect 50498 51652 50522 51654
rect 50282 51632 50578 51652
rect 50282 50620 50578 50640
rect 50338 50618 50362 50620
rect 50418 50618 50442 50620
rect 50498 50618 50522 50620
rect 50360 50566 50362 50618
rect 50424 50566 50436 50618
rect 50498 50566 50500 50618
rect 50338 50564 50362 50566
rect 50418 50564 50442 50566
rect 50498 50564 50522 50566
rect 50282 50544 50578 50564
rect 50282 49532 50578 49552
rect 50338 49530 50362 49532
rect 50418 49530 50442 49532
rect 50498 49530 50522 49532
rect 50360 49478 50362 49530
rect 50424 49478 50436 49530
rect 50498 49478 50500 49530
rect 50338 49476 50362 49478
rect 50418 49476 50442 49478
rect 50498 49476 50522 49478
rect 50282 49456 50578 49476
rect 50282 48444 50578 48464
rect 50338 48442 50362 48444
rect 50418 48442 50442 48444
rect 50498 48442 50522 48444
rect 50360 48390 50362 48442
rect 50424 48390 50436 48442
rect 50498 48390 50500 48442
rect 50338 48388 50362 48390
rect 50418 48388 50442 48390
rect 50498 48388 50522 48390
rect 50282 48368 50578 48388
rect 51166 48278 51194 53094
rect 51154 48272 51206 48278
rect 51154 48214 51206 48220
rect 51246 48272 51298 48278
rect 51246 48214 51298 48220
rect 50282 47356 50578 47376
rect 50338 47354 50362 47356
rect 50418 47354 50442 47356
rect 50498 47354 50522 47356
rect 50360 47302 50362 47354
rect 50424 47302 50436 47354
rect 50498 47302 50500 47354
rect 50338 47300 50362 47302
rect 50418 47300 50442 47302
rect 50498 47300 50522 47302
rect 50282 47280 50578 47300
rect 50282 46268 50578 46288
rect 50338 46266 50362 46268
rect 50418 46266 50442 46268
rect 50498 46266 50522 46268
rect 50360 46214 50362 46266
rect 50424 46214 50436 46266
rect 50498 46214 50500 46266
rect 50338 46212 50362 46214
rect 50418 46212 50442 46214
rect 50498 46212 50522 46214
rect 50282 46192 50578 46212
rect 50282 45180 50578 45200
rect 50338 45178 50362 45180
rect 50418 45178 50442 45180
rect 50498 45178 50522 45180
rect 50360 45126 50362 45178
rect 50424 45126 50436 45178
rect 50498 45126 50500 45178
rect 50338 45124 50362 45126
rect 50418 45124 50442 45126
rect 50498 45124 50522 45126
rect 50282 45104 50578 45124
rect 50282 44092 50578 44112
rect 50338 44090 50362 44092
rect 50418 44090 50442 44092
rect 50498 44090 50522 44092
rect 50360 44038 50362 44090
rect 50424 44038 50436 44090
rect 50498 44038 50500 44090
rect 50338 44036 50362 44038
rect 50418 44036 50442 44038
rect 50498 44036 50522 44038
rect 50282 44016 50578 44036
rect 50970 43784 51022 43790
rect 51062 43784 51114 43790
rect 51022 43732 51062 43738
rect 50970 43726 51114 43732
rect 50982 43710 51102 43726
rect 51258 43330 51286 48214
rect 51074 43302 51286 43330
rect 50282 43004 50578 43024
rect 50338 43002 50362 43004
rect 50418 43002 50442 43004
rect 50498 43002 50522 43004
rect 50360 42950 50362 43002
rect 50424 42950 50436 43002
rect 50498 42950 50500 43002
rect 50338 42948 50362 42950
rect 50418 42948 50442 42950
rect 50498 42948 50522 42950
rect 50282 42928 50578 42948
rect 50282 41916 50578 41936
rect 50338 41914 50362 41916
rect 50418 41914 50442 41916
rect 50498 41914 50522 41916
rect 50360 41862 50362 41914
rect 50424 41862 50436 41914
rect 50498 41862 50500 41914
rect 50338 41860 50362 41862
rect 50418 41860 50442 41862
rect 50498 41860 50522 41862
rect 50282 41840 50578 41860
rect 50282 40828 50578 40848
rect 50338 40826 50362 40828
rect 50418 40826 50442 40828
rect 50498 40826 50522 40828
rect 50360 40774 50362 40826
rect 50424 40774 50436 40826
rect 50498 40774 50500 40826
rect 50338 40772 50362 40774
rect 50418 40772 50442 40774
rect 50498 40772 50522 40774
rect 50282 40752 50578 40772
rect 50970 40384 51022 40390
rect 50970 40326 51022 40332
rect 50282 39740 50578 39760
rect 50338 39738 50362 39740
rect 50418 39738 50442 39740
rect 50498 39738 50522 39740
rect 50360 39686 50362 39738
rect 50424 39686 50436 39738
rect 50498 39686 50500 39738
rect 50338 39684 50362 39686
rect 50418 39684 50442 39686
rect 50498 39684 50522 39686
rect 50282 39664 50578 39684
rect 50282 38652 50578 38672
rect 50338 38650 50362 38652
rect 50418 38650 50442 38652
rect 50498 38650 50522 38652
rect 50360 38598 50362 38650
rect 50424 38598 50436 38650
rect 50498 38598 50500 38650
rect 50338 38596 50362 38598
rect 50418 38596 50442 38598
rect 50498 38596 50522 38598
rect 50282 38576 50578 38596
rect 50282 37564 50578 37584
rect 50338 37562 50362 37564
rect 50418 37562 50442 37564
rect 50498 37562 50522 37564
rect 50360 37510 50362 37562
rect 50424 37510 50436 37562
rect 50498 37510 50500 37562
rect 50338 37508 50362 37510
rect 50418 37508 50442 37510
rect 50498 37508 50522 37510
rect 50282 37488 50578 37508
rect 50282 36476 50578 36496
rect 50338 36474 50362 36476
rect 50418 36474 50442 36476
rect 50498 36474 50522 36476
rect 50360 36422 50362 36474
rect 50424 36422 50436 36474
rect 50498 36422 50500 36474
rect 50338 36420 50362 36422
rect 50418 36420 50442 36422
rect 50498 36420 50522 36422
rect 50282 36400 50578 36420
rect 50282 35388 50578 35408
rect 50338 35386 50362 35388
rect 50418 35386 50442 35388
rect 50498 35386 50522 35388
rect 50360 35334 50362 35386
rect 50424 35334 50436 35386
rect 50498 35334 50500 35386
rect 50338 35332 50362 35334
rect 50418 35332 50442 35334
rect 50498 35332 50522 35334
rect 50282 35312 50578 35332
rect 50282 34300 50578 34320
rect 50338 34298 50362 34300
rect 50418 34298 50442 34300
rect 50498 34298 50522 34300
rect 50360 34246 50362 34298
rect 50424 34246 50436 34298
rect 50498 34246 50500 34298
rect 50338 34244 50362 34246
rect 50418 34244 50442 34246
rect 50498 34244 50522 34246
rect 50282 34224 50578 34244
rect 50282 33212 50578 33232
rect 50338 33210 50362 33212
rect 50418 33210 50442 33212
rect 50498 33210 50522 33212
rect 50360 33158 50362 33210
rect 50424 33158 50436 33210
rect 50498 33158 50500 33210
rect 50338 33156 50362 33158
rect 50418 33156 50442 33158
rect 50498 33156 50522 33158
rect 50282 33136 50578 33156
rect 50282 32124 50578 32144
rect 50338 32122 50362 32124
rect 50418 32122 50442 32124
rect 50498 32122 50522 32124
rect 50360 32070 50362 32122
rect 50424 32070 50436 32122
rect 50498 32070 50500 32122
rect 50338 32068 50362 32070
rect 50418 32068 50442 32070
rect 50498 32068 50522 32070
rect 50282 32048 50578 32068
rect 50282 31036 50578 31056
rect 50338 31034 50362 31036
rect 50418 31034 50442 31036
rect 50498 31034 50522 31036
rect 50360 30982 50362 31034
rect 50424 30982 50436 31034
rect 50498 30982 50500 31034
rect 50338 30980 50362 30982
rect 50418 30980 50442 30982
rect 50498 30980 50522 30982
rect 50282 30960 50578 30980
rect 50282 29948 50578 29968
rect 50338 29946 50362 29948
rect 50418 29946 50442 29948
rect 50498 29946 50522 29948
rect 50360 29894 50362 29946
rect 50424 29894 50436 29946
rect 50498 29894 50500 29946
rect 50338 29892 50362 29894
rect 50418 29892 50442 29894
rect 50498 29892 50522 29894
rect 50282 29872 50578 29892
rect 50282 28860 50578 28880
rect 50338 28858 50362 28860
rect 50418 28858 50442 28860
rect 50498 28858 50522 28860
rect 50360 28806 50362 28858
rect 50424 28806 50436 28858
rect 50498 28806 50500 28858
rect 50338 28804 50362 28806
rect 50418 28804 50442 28806
rect 50498 28804 50522 28806
rect 50282 28784 50578 28804
rect 50282 27772 50578 27792
rect 50338 27770 50362 27772
rect 50418 27770 50442 27772
rect 50498 27770 50522 27772
rect 50360 27718 50362 27770
rect 50424 27718 50436 27770
rect 50498 27718 50500 27770
rect 50338 27716 50362 27718
rect 50418 27716 50442 27718
rect 50498 27716 50522 27718
rect 50282 27696 50578 27716
rect 50282 26684 50578 26704
rect 50338 26682 50362 26684
rect 50418 26682 50442 26684
rect 50498 26682 50522 26684
rect 50360 26630 50362 26682
rect 50424 26630 50436 26682
rect 50498 26630 50500 26682
rect 50338 26628 50362 26630
rect 50418 26628 50442 26630
rect 50498 26628 50522 26630
rect 50282 26608 50578 26628
rect 50282 25596 50578 25616
rect 50338 25594 50362 25596
rect 50418 25594 50442 25596
rect 50498 25594 50522 25596
rect 50360 25542 50362 25594
rect 50424 25542 50436 25594
rect 50498 25542 50500 25594
rect 50338 25540 50362 25542
rect 50418 25540 50442 25542
rect 50498 25540 50522 25542
rect 50282 25520 50578 25540
rect 50282 24508 50578 24528
rect 50338 24506 50362 24508
rect 50418 24506 50442 24508
rect 50498 24506 50522 24508
rect 50360 24454 50362 24506
rect 50424 24454 50436 24506
rect 50498 24454 50500 24506
rect 50338 24452 50362 24454
rect 50418 24452 50442 24454
rect 50498 24452 50522 24454
rect 50282 24432 50578 24452
rect 50282 23420 50578 23440
rect 50338 23418 50362 23420
rect 50418 23418 50442 23420
rect 50498 23418 50522 23420
rect 50360 23366 50362 23418
rect 50424 23366 50436 23418
rect 50498 23366 50500 23418
rect 50338 23364 50362 23366
rect 50418 23364 50442 23366
rect 50498 23364 50522 23366
rect 50282 23344 50578 23364
rect 50282 22332 50578 22352
rect 50338 22330 50362 22332
rect 50418 22330 50442 22332
rect 50498 22330 50522 22332
rect 50360 22278 50362 22330
rect 50424 22278 50436 22330
rect 50498 22278 50500 22330
rect 50338 22276 50362 22278
rect 50418 22276 50442 22278
rect 50498 22276 50522 22278
rect 50282 22256 50578 22276
rect 50602 21956 50654 21962
rect 50602 21898 50654 21904
rect 50282 21244 50578 21264
rect 50338 21242 50362 21244
rect 50418 21242 50442 21244
rect 50498 21242 50522 21244
rect 50360 21190 50362 21242
rect 50424 21190 50436 21242
rect 50498 21190 50500 21242
rect 50338 21188 50362 21190
rect 50418 21188 50442 21190
rect 50498 21188 50522 21190
rect 50282 21168 50578 21188
rect 50282 20156 50578 20176
rect 50338 20154 50362 20156
rect 50418 20154 50442 20156
rect 50498 20154 50522 20156
rect 50360 20102 50362 20154
rect 50424 20102 50436 20154
rect 50498 20102 50500 20154
rect 50338 20100 50362 20102
rect 50418 20100 50442 20102
rect 50498 20100 50522 20102
rect 50282 20080 50578 20100
rect 50282 19068 50578 19088
rect 50338 19066 50362 19068
rect 50418 19066 50442 19068
rect 50498 19066 50522 19068
rect 50360 19014 50362 19066
rect 50424 19014 50436 19066
rect 50498 19014 50500 19066
rect 50338 19012 50362 19014
rect 50418 19012 50442 19014
rect 50498 19012 50522 19014
rect 50282 18992 50578 19012
rect 50282 17980 50578 18000
rect 50338 17978 50362 17980
rect 50418 17978 50442 17980
rect 50498 17978 50522 17980
rect 50360 17926 50362 17978
rect 50424 17926 50436 17978
rect 50498 17926 50500 17978
rect 50338 17924 50362 17926
rect 50418 17924 50442 17926
rect 50498 17924 50522 17926
rect 50282 17904 50578 17924
rect 50282 16892 50578 16912
rect 50338 16890 50362 16892
rect 50418 16890 50442 16892
rect 50498 16890 50522 16892
rect 50360 16838 50362 16890
rect 50424 16838 50436 16890
rect 50498 16838 50500 16890
rect 50338 16836 50362 16838
rect 50418 16836 50442 16838
rect 50498 16836 50522 16838
rect 50282 16816 50578 16836
rect 50282 15804 50578 15824
rect 50338 15802 50362 15804
rect 50418 15802 50442 15804
rect 50498 15802 50522 15804
rect 50360 15750 50362 15802
rect 50424 15750 50436 15802
rect 50498 15750 50500 15802
rect 50338 15748 50362 15750
rect 50418 15748 50442 15750
rect 50498 15748 50522 15750
rect 50282 15728 50578 15748
rect 50282 14716 50578 14736
rect 50338 14714 50362 14716
rect 50418 14714 50442 14716
rect 50498 14714 50522 14716
rect 50360 14662 50362 14714
rect 50424 14662 50436 14714
rect 50498 14662 50500 14714
rect 50338 14660 50362 14662
rect 50418 14660 50442 14662
rect 50498 14660 50522 14662
rect 50282 14640 50578 14660
rect 49866 13796 49918 13802
rect 49866 13738 49918 13744
rect 50282 13628 50578 13648
rect 50338 13626 50362 13628
rect 50418 13626 50442 13628
rect 50498 13626 50522 13628
rect 50360 13574 50362 13626
rect 50424 13574 50436 13626
rect 50498 13574 50500 13626
rect 50338 13572 50362 13574
rect 50418 13572 50442 13574
rect 50498 13572 50522 13574
rect 50282 13552 50578 13572
rect 50282 12540 50578 12560
rect 50338 12538 50362 12540
rect 50418 12538 50442 12540
rect 50498 12538 50522 12540
rect 50360 12486 50362 12538
rect 50424 12486 50436 12538
rect 50498 12486 50500 12538
rect 50338 12484 50362 12486
rect 50418 12484 50442 12486
rect 50498 12484 50522 12486
rect 50282 12464 50578 12484
rect 50282 11452 50578 11472
rect 50338 11450 50362 11452
rect 50418 11450 50442 11452
rect 50498 11450 50522 11452
rect 50360 11398 50362 11450
rect 50424 11398 50436 11450
rect 50498 11398 50500 11450
rect 50338 11396 50362 11398
rect 50418 11396 50442 11398
rect 50498 11396 50522 11398
rect 50282 11376 50578 11396
rect 50282 10364 50578 10384
rect 50338 10362 50362 10364
rect 50418 10362 50442 10364
rect 50498 10362 50522 10364
rect 50360 10310 50362 10362
rect 50424 10310 50436 10362
rect 50498 10310 50500 10362
rect 50338 10308 50362 10310
rect 50418 10308 50442 10310
rect 50498 10308 50522 10310
rect 50282 10288 50578 10308
rect 50142 9920 50194 9926
rect 50142 9862 50194 9868
rect 49774 4004 49826 4010
rect 49774 3946 49826 3952
rect 49682 3120 49734 3126
rect 49682 3062 49734 3068
rect 49694 2854 49722 3062
rect 49682 2848 49734 2854
rect 49682 2790 49734 2796
rect 49418 870 49630 898
rect 49418 800 49446 870
rect 49786 800 49814 3946
rect 49958 3664 50010 3670
rect 49958 3606 50010 3612
rect 49970 1426 49998 3606
rect 50154 3602 50182 9862
rect 50282 9276 50578 9296
rect 50338 9274 50362 9276
rect 50418 9274 50442 9276
rect 50498 9274 50522 9276
rect 50360 9222 50362 9274
rect 50424 9222 50436 9274
rect 50498 9222 50500 9274
rect 50338 9220 50362 9222
rect 50418 9220 50442 9222
rect 50498 9220 50522 9222
rect 50282 9200 50578 9220
rect 50282 8188 50578 8208
rect 50338 8186 50362 8188
rect 50418 8186 50442 8188
rect 50498 8186 50522 8188
rect 50360 8134 50362 8186
rect 50424 8134 50436 8186
rect 50498 8134 50500 8186
rect 50338 8132 50362 8134
rect 50418 8132 50442 8134
rect 50498 8132 50522 8134
rect 50282 8112 50578 8132
rect 50282 7100 50578 7120
rect 50338 7098 50362 7100
rect 50418 7098 50442 7100
rect 50498 7098 50522 7100
rect 50360 7046 50362 7098
rect 50424 7046 50436 7098
rect 50498 7046 50500 7098
rect 50338 7044 50362 7046
rect 50418 7044 50442 7046
rect 50498 7044 50522 7046
rect 50282 7024 50578 7044
rect 50282 6012 50578 6032
rect 50338 6010 50362 6012
rect 50418 6010 50442 6012
rect 50498 6010 50522 6012
rect 50360 5958 50362 6010
rect 50424 5958 50436 6010
rect 50498 5958 50500 6010
rect 50338 5956 50362 5958
rect 50418 5956 50442 5958
rect 50498 5956 50522 5958
rect 50282 5936 50578 5956
rect 50282 4924 50578 4944
rect 50338 4922 50362 4924
rect 50418 4922 50442 4924
rect 50498 4922 50522 4924
rect 50360 4870 50362 4922
rect 50424 4870 50436 4922
rect 50498 4870 50500 4922
rect 50338 4868 50362 4870
rect 50418 4868 50442 4870
rect 50498 4868 50522 4870
rect 50282 4848 50578 4868
rect 50282 3836 50578 3856
rect 50338 3834 50362 3836
rect 50418 3834 50442 3836
rect 50498 3834 50522 3836
rect 50360 3782 50362 3834
rect 50424 3782 50436 3834
rect 50498 3782 50500 3834
rect 50338 3780 50362 3782
rect 50418 3780 50442 3782
rect 50498 3780 50522 3782
rect 50282 3760 50578 3780
rect 50142 3596 50194 3602
rect 50142 3538 50194 3544
rect 50614 3194 50642 21898
rect 50694 15428 50746 15434
rect 50694 15370 50746 15376
rect 50142 3188 50194 3194
rect 50142 3130 50194 3136
rect 50602 3188 50654 3194
rect 50602 3130 50654 3136
rect 50050 2848 50102 2854
rect 50050 2790 50102 2796
rect 50062 2378 50090 2790
rect 50050 2372 50102 2378
rect 50050 2314 50102 2320
rect 49958 1420 50010 1426
rect 49958 1362 50010 1368
rect 50154 800 50182 3130
rect 50706 3126 50734 15370
rect 50786 4140 50838 4146
rect 50786 4082 50838 4088
rect 50510 3120 50562 3126
rect 50694 3120 50746 3126
rect 50562 3068 50642 3074
rect 50510 3062 50642 3068
rect 50694 3062 50746 3068
rect 50522 3046 50642 3062
rect 50282 2748 50578 2768
rect 50338 2746 50362 2748
rect 50418 2746 50442 2748
rect 50498 2746 50522 2748
rect 50360 2694 50362 2746
rect 50424 2694 50436 2746
rect 50498 2694 50500 2746
rect 50338 2692 50362 2694
rect 50418 2692 50442 2694
rect 50498 2692 50522 2694
rect 50282 2672 50578 2692
rect 50614 1442 50642 3046
rect 50798 2922 50826 4082
rect 50982 4010 51010 40326
rect 51074 31770 51102 43302
rect 51074 31742 51286 31770
rect 51258 19378 51286 31742
rect 51062 19372 51114 19378
rect 51062 19314 51114 19320
rect 51246 19372 51298 19378
rect 51246 19314 51298 19320
rect 51074 16454 51102 19314
rect 51706 18216 51758 18222
rect 51706 18158 51758 18164
rect 51062 16448 51114 16454
rect 51062 16390 51114 16396
rect 51614 4072 51666 4078
rect 51614 4014 51666 4020
rect 50970 4004 51022 4010
rect 50970 3946 51022 3952
rect 51246 3664 51298 3670
rect 51246 3606 51298 3612
rect 50786 2916 50838 2922
rect 50786 2858 50838 2864
rect 50522 1414 50642 1442
rect 50878 1420 50930 1426
rect 50522 800 50550 1414
rect 50878 1362 50930 1368
rect 50890 800 50918 1362
rect 51258 800 51286 3606
rect 51626 800 51654 4014
rect 51718 3738 51746 18158
rect 52350 14272 52402 14278
rect 52350 14214 52402 14220
rect 51798 12776 51850 12782
rect 51798 12718 51850 12724
rect 51810 4146 51838 12718
rect 51798 4140 51850 4146
rect 51798 4082 51850 4088
rect 51706 3732 51758 3738
rect 51706 3674 51758 3680
rect 51982 3052 52034 3058
rect 51982 2994 52034 3000
rect 51994 800 52022 2994
rect 52362 800 52390 14214
rect 52454 898 52482 55558
rect 55110 46504 55162 46510
rect 55110 46446 55162 46452
rect 54190 4140 54242 4146
rect 54190 4082 54242 4088
rect 53822 3528 53874 3534
rect 53822 3470 53874 3476
rect 53454 2916 53506 2922
rect 53454 2858 53506 2864
rect 53086 2576 53138 2582
rect 53086 2518 53138 2524
rect 52454 870 52758 898
rect 52730 800 52758 870
rect 53098 800 53126 2518
rect 53466 800 53494 2858
rect 53834 800 53862 3470
rect 54202 800 54230 4082
rect 54926 3596 54978 3602
rect 54926 3538 54978 3544
rect 54558 3052 54610 3058
rect 54558 2994 54610 3000
rect 54570 800 54598 2994
rect 54938 800 54966 3538
rect 55122 3058 55150 46446
rect 55214 17746 55242 59078
rect 55950 56166 55978 59200
rect 55938 56160 55990 56166
rect 55938 56102 55990 56108
rect 56410 55865 56438 59200
rect 56962 58041 56990 59200
rect 56764 58032 56820 58041
rect 56764 57967 56820 57976
rect 56948 58032 57004 58041
rect 56948 57967 57004 57976
rect 56778 57934 56806 57967
rect 56766 57928 56818 57934
rect 56766 57870 56818 57876
rect 56858 57928 56910 57934
rect 56858 57870 56910 57876
rect 56396 55856 56452 55865
rect 56396 55791 56452 55800
rect 56870 38865 56898 57870
rect 57514 56302 57542 59200
rect 57502 56296 57554 56302
rect 57502 56238 57554 56244
rect 58066 55962 58094 59200
rect 58054 55956 58106 55962
rect 58054 55898 58106 55904
rect 59078 55894 59106 59200
rect 59066 55888 59118 55894
rect 59066 55830 59118 55836
rect 59630 55826 59658 59200
rect 59618 55820 59670 55826
rect 59618 55762 59670 55768
rect 56856 38856 56912 38865
rect 56856 38791 56912 38800
rect 56764 38720 56820 38729
rect 56764 38655 56820 38664
rect 55662 35624 55714 35630
rect 55662 35566 55714 35572
rect 55202 17740 55254 17746
rect 55202 17682 55254 17688
rect 55674 4706 55702 35566
rect 56778 33810 56806 38655
rect 56594 33782 56806 33810
rect 56594 24206 56622 33782
rect 56582 24200 56634 24206
rect 56582 24142 56634 24148
rect 56766 24200 56818 24206
rect 56766 24142 56818 24148
rect 56778 17814 56806 24142
rect 56766 17808 56818 17814
rect 56766 17750 56818 17756
rect 59710 11688 59762 11694
rect 59710 11630 59762 11636
rect 58606 11620 58658 11626
rect 58606 11562 58658 11568
rect 57132 9616 57188 9625
rect 57132 9551 57188 9560
rect 55674 4678 56070 4706
rect 55294 3392 55346 3398
rect 55294 3334 55346 3340
rect 55110 3052 55162 3058
rect 55110 2994 55162 3000
rect 55306 800 55334 3334
rect 55660 2952 55716 2961
rect 55660 2887 55716 2896
rect 55674 800 55702 2887
rect 56042 800 56070 4678
rect 56766 3936 56818 3942
rect 56766 3878 56818 3884
rect 56398 2984 56450 2990
rect 56398 2926 56450 2932
rect 56410 800 56438 2926
rect 56778 800 56806 3878
rect 57146 800 57174 9551
rect 57502 3664 57554 3670
rect 57502 3606 57554 3612
rect 57514 800 57542 3606
rect 58238 3120 58290 3126
rect 58238 3062 58290 3068
rect 57870 2848 57922 2854
rect 57870 2790 57922 2796
rect 57882 800 57910 2790
rect 58250 800 58278 3062
rect 58618 800 58646 11562
rect 59342 3732 59394 3738
rect 59342 3674 59394 3680
rect 58974 3188 59026 3194
rect 58974 3130 59026 3136
rect 58986 800 59014 3130
rect 59354 800 59382 3674
rect 59722 800 59750 11630
rect 0 0 56 800
rect 92 0 148 800
rect 184 0 240 800
rect 276 0 332 800
rect 460 0 516 800
rect 552 0 608 800
rect 644 0 700 800
rect 828 0 884 800
rect 920 0 976 800
rect 1012 0 1068 800
rect 1196 0 1252 800
rect 1288 0 1344 800
rect 1380 0 1436 800
rect 1564 0 1620 800
rect 1656 0 1712 800
rect 1748 0 1804 800
rect 1932 0 1988 800
rect 2024 0 2080 800
rect 2116 0 2172 800
rect 2300 0 2356 800
rect 2392 0 2448 800
rect 2484 0 2540 800
rect 2668 0 2724 800
rect 2760 0 2816 800
rect 2852 0 2908 800
rect 3036 0 3092 800
rect 3128 0 3184 800
rect 3220 0 3276 800
rect 3404 0 3460 800
rect 3496 0 3552 800
rect 3588 0 3644 800
rect 3772 0 3828 800
rect 3864 0 3920 800
rect 3956 0 4012 800
rect 4140 0 4196 800
rect 4232 0 4288 800
rect 4324 0 4380 800
rect 4508 0 4564 800
rect 4600 0 4656 800
rect 4692 0 4748 800
rect 4876 0 4932 800
rect 4968 0 5024 800
rect 5060 0 5116 800
rect 5244 0 5300 800
rect 5336 0 5392 800
rect 5428 0 5484 800
rect 5612 0 5668 800
rect 5704 0 5760 800
rect 5796 0 5852 800
rect 5980 0 6036 800
rect 6072 0 6128 800
rect 6164 0 6220 800
rect 6348 0 6404 800
rect 6440 0 6496 800
rect 6532 0 6588 800
rect 6716 0 6772 800
rect 6808 0 6864 800
rect 6900 0 6956 800
rect 7084 0 7140 800
rect 7176 0 7232 800
rect 7268 0 7324 800
rect 7452 0 7508 800
rect 7544 0 7600 800
rect 7636 0 7692 800
rect 7820 0 7876 800
rect 7912 0 7968 800
rect 8004 0 8060 800
rect 8188 0 8244 800
rect 8280 0 8336 800
rect 8372 0 8428 800
rect 8556 0 8612 800
rect 8648 0 8704 800
rect 8740 0 8796 800
rect 8924 0 8980 800
rect 9016 0 9072 800
rect 9108 0 9164 800
rect 9292 0 9348 800
rect 9384 0 9440 800
rect 9476 0 9532 800
rect 9660 0 9716 800
rect 9752 0 9808 800
rect 9844 0 9900 800
rect 10028 0 10084 800
rect 10120 0 10176 800
rect 10212 0 10268 800
rect 10396 0 10452 800
rect 10488 0 10544 800
rect 10580 0 10636 800
rect 10764 0 10820 800
rect 10856 0 10912 800
rect 10948 0 11004 800
rect 11132 0 11188 800
rect 11224 0 11280 800
rect 11316 0 11372 800
rect 11500 0 11556 800
rect 11592 0 11648 800
rect 11684 0 11740 800
rect 11868 0 11924 800
rect 11960 0 12016 800
rect 12052 0 12108 800
rect 12236 0 12292 800
rect 12328 0 12384 800
rect 12420 0 12476 800
rect 12604 0 12660 800
rect 12696 0 12752 800
rect 12788 0 12844 800
rect 12972 0 13028 800
rect 13064 0 13120 800
rect 13156 0 13212 800
rect 13340 0 13396 800
rect 13432 0 13488 800
rect 13524 0 13580 800
rect 13708 0 13764 800
rect 13800 0 13856 800
rect 13892 0 13948 800
rect 14076 0 14132 800
rect 14168 0 14224 800
rect 14260 0 14316 800
rect 14444 0 14500 800
rect 14536 0 14592 800
rect 14628 0 14684 800
rect 14812 0 14868 800
rect 14904 0 14960 800
rect 14996 0 15052 800
rect 15088 0 15144 800
rect 15272 0 15328 800
rect 15364 0 15420 800
rect 15456 0 15512 800
rect 15640 0 15696 800
rect 15732 0 15788 800
rect 15824 0 15880 800
rect 16008 0 16064 800
rect 16100 0 16156 800
rect 16192 0 16248 800
rect 16376 0 16432 800
rect 16468 0 16524 800
rect 16560 0 16616 800
rect 16744 0 16800 800
rect 16836 0 16892 800
rect 16928 0 16984 800
rect 17112 0 17168 800
rect 17204 0 17260 800
rect 17296 0 17352 800
rect 17480 0 17536 800
rect 17572 0 17628 800
rect 17664 0 17720 800
rect 17848 0 17904 800
rect 17940 0 17996 800
rect 18032 0 18088 800
rect 18216 0 18272 800
rect 18308 0 18364 800
rect 18400 0 18456 800
rect 18584 0 18640 800
rect 18676 0 18732 800
rect 18768 0 18824 800
rect 18952 0 19008 800
rect 19044 0 19100 800
rect 19136 0 19192 800
rect 19320 0 19376 800
rect 19412 0 19468 800
rect 19504 0 19560 800
rect 19688 0 19744 800
rect 19780 0 19836 800
rect 19872 0 19928 800
rect 20056 0 20112 800
rect 20148 0 20204 800
rect 20240 0 20296 800
rect 20424 0 20480 800
rect 20516 0 20572 800
rect 20608 0 20664 800
rect 20792 0 20848 800
rect 20884 0 20940 800
rect 20976 0 21032 800
rect 21160 0 21216 800
rect 21252 0 21308 800
rect 21344 0 21400 800
rect 21528 0 21584 800
rect 21620 0 21676 800
rect 21712 0 21768 800
rect 21896 0 21952 800
rect 21988 0 22044 800
rect 22080 0 22136 800
rect 22264 0 22320 800
rect 22356 0 22412 800
rect 22448 0 22504 800
rect 22632 0 22688 800
rect 22724 0 22780 800
rect 22816 0 22872 800
rect 23000 0 23056 800
rect 23092 0 23148 800
rect 23184 0 23240 800
rect 23368 0 23424 800
rect 23460 0 23516 800
rect 23552 0 23608 800
rect 23736 0 23792 800
rect 23828 0 23884 800
rect 23920 0 23976 800
rect 24104 0 24160 800
rect 24196 0 24252 800
rect 24288 0 24344 800
rect 24472 0 24528 800
rect 24564 0 24620 800
rect 24656 0 24712 800
rect 24840 0 24896 800
rect 24932 0 24988 800
rect 25024 0 25080 800
rect 25208 0 25264 800
rect 25300 0 25356 800
rect 25392 0 25448 800
rect 25576 0 25632 800
rect 25668 0 25724 800
rect 25760 0 25816 800
rect 25944 0 26000 800
rect 26036 0 26092 800
rect 26128 0 26184 800
rect 26312 0 26368 800
rect 26404 0 26460 800
rect 26496 0 26552 800
rect 26680 0 26736 800
rect 26772 0 26828 800
rect 26864 0 26920 800
rect 27048 0 27104 800
rect 27140 0 27196 800
rect 27232 0 27288 800
rect 27416 0 27472 800
rect 27508 0 27564 800
rect 27600 0 27656 800
rect 27784 0 27840 800
rect 27876 0 27932 800
rect 27968 0 28024 800
rect 28152 0 28208 800
rect 28244 0 28300 800
rect 28336 0 28392 800
rect 28520 0 28576 800
rect 28612 0 28668 800
rect 28704 0 28760 800
rect 28888 0 28944 800
rect 28980 0 29036 800
rect 29072 0 29128 800
rect 29256 0 29312 800
rect 29348 0 29404 800
rect 29440 0 29496 800
rect 29624 0 29680 800
rect 29716 0 29772 800
rect 29808 0 29864 800
rect 29992 0 30048 800
rect 30084 0 30140 800
rect 30176 0 30232 800
rect 30268 0 30324 800
rect 30452 0 30508 800
rect 30544 0 30600 800
rect 30636 0 30692 800
rect 30820 0 30876 800
rect 30912 0 30968 800
rect 31004 0 31060 800
rect 31188 0 31244 800
rect 31280 0 31336 800
rect 31372 0 31428 800
rect 31556 0 31612 800
rect 31648 0 31704 800
rect 31740 0 31796 800
rect 31924 0 31980 800
rect 32016 0 32072 800
rect 32108 0 32164 800
rect 32292 0 32348 800
rect 32384 0 32440 800
rect 32476 0 32532 800
rect 32660 0 32716 800
rect 32752 0 32808 800
rect 32844 0 32900 800
rect 33028 0 33084 800
rect 33120 0 33176 800
rect 33212 0 33268 800
rect 33396 0 33452 800
rect 33488 0 33544 800
rect 33580 0 33636 800
rect 33764 0 33820 800
rect 33856 0 33912 800
rect 33948 0 34004 800
rect 34132 0 34188 800
rect 34224 0 34280 800
rect 34316 0 34372 800
rect 34500 0 34556 800
rect 34592 0 34648 800
rect 34684 0 34740 800
rect 34868 0 34924 800
rect 34960 0 35016 800
rect 35052 0 35108 800
rect 35236 0 35292 800
rect 35328 0 35384 800
rect 35420 0 35476 800
rect 35604 0 35660 800
rect 35696 0 35752 800
rect 35788 0 35844 800
rect 35972 0 36028 800
rect 36064 0 36120 800
rect 36156 0 36212 800
rect 36340 0 36396 800
rect 36432 0 36488 800
rect 36524 0 36580 800
rect 36708 0 36764 800
rect 36800 0 36856 800
rect 36892 0 36948 800
rect 37076 0 37132 800
rect 37168 0 37224 800
rect 37260 0 37316 800
rect 37444 0 37500 800
rect 37536 0 37592 800
rect 37628 0 37684 800
rect 37812 0 37868 800
rect 37904 0 37960 800
rect 37996 0 38052 800
rect 38180 0 38236 800
rect 38272 0 38328 800
rect 38364 0 38420 800
rect 38548 0 38604 800
rect 38640 0 38696 800
rect 38732 0 38788 800
rect 38916 0 38972 800
rect 39008 0 39064 800
rect 39100 0 39156 800
rect 39284 0 39340 800
rect 39376 0 39432 800
rect 39468 0 39524 800
rect 39652 0 39708 800
rect 39744 0 39800 800
rect 39836 0 39892 800
rect 40020 0 40076 800
rect 40112 0 40168 800
rect 40204 0 40260 800
rect 40388 0 40444 800
rect 40480 0 40536 800
rect 40572 0 40628 800
rect 40756 0 40812 800
rect 40848 0 40904 800
rect 40940 0 40996 800
rect 41124 0 41180 800
rect 41216 0 41272 800
rect 41308 0 41364 800
rect 41492 0 41548 800
rect 41584 0 41640 800
rect 41676 0 41732 800
rect 41860 0 41916 800
rect 41952 0 42008 800
rect 42044 0 42100 800
rect 42228 0 42284 800
rect 42320 0 42376 800
rect 42412 0 42468 800
rect 42596 0 42652 800
rect 42688 0 42744 800
rect 42780 0 42836 800
rect 42964 0 43020 800
rect 43056 0 43112 800
rect 43148 0 43204 800
rect 43332 0 43388 800
rect 43424 0 43480 800
rect 43516 0 43572 800
rect 43700 0 43756 800
rect 43792 0 43848 800
rect 43884 0 43940 800
rect 44068 0 44124 800
rect 44160 0 44216 800
rect 44252 0 44308 800
rect 44436 0 44492 800
rect 44528 0 44584 800
rect 44620 0 44676 800
rect 44804 0 44860 800
rect 44896 0 44952 800
rect 44988 0 45044 800
rect 45080 0 45136 800
rect 45264 0 45320 800
rect 45356 0 45412 800
rect 45448 0 45504 800
rect 45632 0 45688 800
rect 45724 0 45780 800
rect 45816 0 45872 800
rect 46000 0 46056 800
rect 46092 0 46148 800
rect 46184 0 46240 800
rect 46368 0 46424 800
rect 46460 0 46516 800
rect 46552 0 46608 800
rect 46736 0 46792 800
rect 46828 0 46884 800
rect 46920 0 46976 800
rect 47104 0 47160 800
rect 47196 0 47252 800
rect 47288 0 47344 800
rect 47472 0 47528 800
rect 47564 0 47620 800
rect 47656 0 47712 800
rect 47840 0 47896 800
rect 47932 0 47988 800
rect 48024 0 48080 800
rect 48208 0 48264 800
rect 48300 0 48356 800
rect 48392 0 48448 800
rect 48576 0 48632 800
rect 48668 0 48724 800
rect 48760 0 48816 800
rect 48944 0 49000 800
rect 49036 0 49092 800
rect 49128 0 49184 800
rect 49312 0 49368 800
rect 49404 0 49460 800
rect 49496 0 49552 800
rect 49680 0 49736 800
rect 49772 0 49828 800
rect 49864 0 49920 800
rect 50048 0 50104 800
rect 50140 0 50196 800
rect 50232 0 50288 800
rect 50416 0 50472 800
rect 50508 0 50564 800
rect 50600 0 50656 800
rect 50784 0 50840 800
rect 50876 0 50932 800
rect 50968 0 51024 800
rect 51152 0 51208 800
rect 51244 0 51300 800
rect 51336 0 51392 800
rect 51520 0 51576 800
rect 51612 0 51668 800
rect 51704 0 51760 800
rect 51888 0 51944 800
rect 51980 0 52036 800
rect 52072 0 52128 800
rect 52256 0 52312 800
rect 52348 0 52404 800
rect 52440 0 52496 800
rect 52624 0 52680 800
rect 52716 0 52772 800
rect 52808 0 52864 800
rect 52992 0 53048 800
rect 53084 0 53140 800
rect 53176 0 53232 800
rect 53360 0 53416 800
rect 53452 0 53508 800
rect 53544 0 53600 800
rect 53728 0 53784 800
rect 53820 0 53876 800
rect 53912 0 53968 800
rect 54096 0 54152 800
rect 54188 0 54244 800
rect 54280 0 54336 800
rect 54464 0 54520 800
rect 54556 0 54612 800
rect 54648 0 54704 800
rect 54832 0 54888 800
rect 54924 0 54980 800
rect 55016 0 55072 800
rect 55200 0 55256 800
rect 55292 0 55348 800
rect 55384 0 55440 800
rect 55568 0 55624 800
rect 55660 0 55716 800
rect 55752 0 55808 800
rect 55936 0 55992 800
rect 56028 0 56084 800
rect 56120 0 56176 800
rect 56304 0 56360 800
rect 56396 0 56452 800
rect 56488 0 56544 800
rect 56672 0 56728 800
rect 56764 0 56820 800
rect 56856 0 56912 800
rect 57040 0 57096 800
rect 57132 0 57188 800
rect 57224 0 57280 800
rect 57408 0 57464 800
rect 57500 0 57556 800
rect 57592 0 57648 800
rect 57776 0 57832 800
rect 57868 0 57924 800
rect 57960 0 58016 800
rect 58144 0 58200 800
rect 58236 0 58292 800
rect 58328 0 58384 800
rect 58512 0 58568 800
rect 58604 0 58660 800
rect 58696 0 58752 800
rect 58880 0 58936 800
rect 58972 0 59028 800
rect 59064 0 59120 800
rect 59248 0 59304 800
rect 59340 0 59396 800
rect 59432 0 59488 800
rect 59616 0 59672 800
rect 59708 0 59764 800
rect 59800 0 59856 800
<< via2 >>
rect 4202 57690 4258 57692
rect 4282 57690 4338 57692
rect 4362 57690 4418 57692
rect 4442 57690 4498 57692
rect 4202 57638 4228 57690
rect 4228 57638 4258 57690
rect 4282 57638 4292 57690
rect 4292 57638 4338 57690
rect 4362 57638 4408 57690
rect 4408 57638 4418 57690
rect 4442 57638 4472 57690
rect 4472 57638 4498 57690
rect 4202 57636 4258 57638
rect 4282 57636 4338 57638
rect 4362 57636 4418 57638
rect 4442 57636 4498 57638
rect 4202 56602 4258 56604
rect 4282 56602 4338 56604
rect 4362 56602 4418 56604
rect 4442 56602 4498 56604
rect 4202 56550 4228 56602
rect 4228 56550 4258 56602
rect 4282 56550 4292 56602
rect 4292 56550 4338 56602
rect 4362 56550 4408 56602
rect 4408 56550 4418 56602
rect 4442 56550 4472 56602
rect 4472 56550 4498 56602
rect 4202 56548 4258 56550
rect 4282 56548 4338 56550
rect 4362 56548 4418 56550
rect 4442 56548 4498 56550
rect 4202 55514 4258 55516
rect 4282 55514 4338 55516
rect 4362 55514 4418 55516
rect 4442 55514 4498 55516
rect 4202 55462 4228 55514
rect 4228 55462 4258 55514
rect 4282 55462 4292 55514
rect 4292 55462 4338 55514
rect 4362 55462 4408 55514
rect 4408 55462 4418 55514
rect 4442 55462 4472 55514
rect 4472 55462 4498 55514
rect 4202 55460 4258 55462
rect 4282 55460 4338 55462
rect 4362 55460 4418 55462
rect 4442 55460 4498 55462
rect 4202 54426 4258 54428
rect 4282 54426 4338 54428
rect 4362 54426 4418 54428
rect 4442 54426 4498 54428
rect 4202 54374 4228 54426
rect 4228 54374 4258 54426
rect 4282 54374 4292 54426
rect 4292 54374 4338 54426
rect 4362 54374 4408 54426
rect 4408 54374 4418 54426
rect 4442 54374 4472 54426
rect 4472 54374 4498 54426
rect 4202 54372 4258 54374
rect 4282 54372 4338 54374
rect 4362 54372 4418 54374
rect 4442 54372 4498 54374
rect 4202 53338 4258 53340
rect 4282 53338 4338 53340
rect 4362 53338 4418 53340
rect 4442 53338 4498 53340
rect 4202 53286 4228 53338
rect 4228 53286 4258 53338
rect 4282 53286 4292 53338
rect 4292 53286 4338 53338
rect 4362 53286 4408 53338
rect 4408 53286 4418 53338
rect 4442 53286 4472 53338
rect 4472 53286 4498 53338
rect 4202 53284 4258 53286
rect 4282 53284 4338 53286
rect 4362 53284 4418 53286
rect 4442 53284 4498 53286
rect 4202 52250 4258 52252
rect 4282 52250 4338 52252
rect 4362 52250 4418 52252
rect 4442 52250 4498 52252
rect 4202 52198 4228 52250
rect 4228 52198 4258 52250
rect 4282 52198 4292 52250
rect 4292 52198 4338 52250
rect 4362 52198 4408 52250
rect 4408 52198 4418 52250
rect 4442 52198 4472 52250
rect 4472 52198 4498 52250
rect 4202 52196 4258 52198
rect 4282 52196 4338 52198
rect 4362 52196 4418 52198
rect 4442 52196 4498 52198
rect 4202 51162 4258 51164
rect 4282 51162 4338 51164
rect 4362 51162 4418 51164
rect 4442 51162 4498 51164
rect 4202 51110 4228 51162
rect 4228 51110 4258 51162
rect 4282 51110 4292 51162
rect 4292 51110 4338 51162
rect 4362 51110 4408 51162
rect 4408 51110 4418 51162
rect 4442 51110 4472 51162
rect 4472 51110 4498 51162
rect 4202 51108 4258 51110
rect 4282 51108 4338 51110
rect 4362 51108 4418 51110
rect 4442 51108 4498 51110
rect 4202 50074 4258 50076
rect 4282 50074 4338 50076
rect 4362 50074 4418 50076
rect 4442 50074 4498 50076
rect 4202 50022 4228 50074
rect 4228 50022 4258 50074
rect 4282 50022 4292 50074
rect 4292 50022 4338 50074
rect 4362 50022 4408 50074
rect 4408 50022 4418 50074
rect 4442 50022 4472 50074
rect 4472 50022 4498 50074
rect 4202 50020 4258 50022
rect 4282 50020 4338 50022
rect 4362 50020 4418 50022
rect 4442 50020 4498 50022
rect 4202 48986 4258 48988
rect 4282 48986 4338 48988
rect 4362 48986 4418 48988
rect 4442 48986 4498 48988
rect 4202 48934 4228 48986
rect 4228 48934 4258 48986
rect 4282 48934 4292 48986
rect 4292 48934 4338 48986
rect 4362 48934 4408 48986
rect 4408 48934 4418 48986
rect 4442 48934 4472 48986
rect 4472 48934 4498 48986
rect 4202 48932 4258 48934
rect 4282 48932 4338 48934
rect 4362 48932 4418 48934
rect 4442 48932 4498 48934
rect 4202 47898 4258 47900
rect 4282 47898 4338 47900
rect 4362 47898 4418 47900
rect 4442 47898 4498 47900
rect 4202 47846 4228 47898
rect 4228 47846 4258 47898
rect 4282 47846 4292 47898
rect 4292 47846 4338 47898
rect 4362 47846 4408 47898
rect 4408 47846 4418 47898
rect 4442 47846 4472 47898
rect 4472 47846 4498 47898
rect 4202 47844 4258 47846
rect 4282 47844 4338 47846
rect 4362 47844 4418 47846
rect 4442 47844 4498 47846
rect 4202 46810 4258 46812
rect 4282 46810 4338 46812
rect 4362 46810 4418 46812
rect 4442 46810 4498 46812
rect 4202 46758 4228 46810
rect 4228 46758 4258 46810
rect 4282 46758 4292 46810
rect 4292 46758 4338 46810
rect 4362 46758 4408 46810
rect 4408 46758 4418 46810
rect 4442 46758 4472 46810
rect 4472 46758 4498 46810
rect 4202 46756 4258 46758
rect 4282 46756 4338 46758
rect 4362 46756 4418 46758
rect 4442 46756 4498 46758
rect 4202 45722 4258 45724
rect 4282 45722 4338 45724
rect 4362 45722 4418 45724
rect 4442 45722 4498 45724
rect 4202 45670 4228 45722
rect 4228 45670 4258 45722
rect 4282 45670 4292 45722
rect 4292 45670 4338 45722
rect 4362 45670 4408 45722
rect 4408 45670 4418 45722
rect 4442 45670 4472 45722
rect 4472 45670 4498 45722
rect 4202 45668 4258 45670
rect 4282 45668 4338 45670
rect 4362 45668 4418 45670
rect 4442 45668 4498 45670
rect 4202 44634 4258 44636
rect 4282 44634 4338 44636
rect 4362 44634 4418 44636
rect 4442 44634 4498 44636
rect 4202 44582 4228 44634
rect 4228 44582 4258 44634
rect 4282 44582 4292 44634
rect 4292 44582 4338 44634
rect 4362 44582 4408 44634
rect 4408 44582 4418 44634
rect 4442 44582 4472 44634
rect 4472 44582 4498 44634
rect 4202 44580 4258 44582
rect 4282 44580 4338 44582
rect 4362 44580 4418 44582
rect 4442 44580 4498 44582
rect 4202 43546 4258 43548
rect 4282 43546 4338 43548
rect 4362 43546 4418 43548
rect 4442 43546 4498 43548
rect 4202 43494 4228 43546
rect 4228 43494 4258 43546
rect 4282 43494 4292 43546
rect 4292 43494 4338 43546
rect 4362 43494 4408 43546
rect 4408 43494 4418 43546
rect 4442 43494 4472 43546
rect 4472 43494 4498 43546
rect 4202 43492 4258 43494
rect 4282 43492 4338 43494
rect 4362 43492 4418 43494
rect 4442 43492 4498 43494
rect 4202 42458 4258 42460
rect 4282 42458 4338 42460
rect 4362 42458 4418 42460
rect 4442 42458 4498 42460
rect 4202 42406 4228 42458
rect 4228 42406 4258 42458
rect 4282 42406 4292 42458
rect 4292 42406 4338 42458
rect 4362 42406 4408 42458
rect 4408 42406 4418 42458
rect 4442 42406 4472 42458
rect 4472 42406 4498 42458
rect 4202 42404 4258 42406
rect 4282 42404 4338 42406
rect 4362 42404 4418 42406
rect 4442 42404 4498 42406
rect 4202 41370 4258 41372
rect 4282 41370 4338 41372
rect 4362 41370 4418 41372
rect 4442 41370 4498 41372
rect 4202 41318 4228 41370
rect 4228 41318 4258 41370
rect 4282 41318 4292 41370
rect 4292 41318 4338 41370
rect 4362 41318 4408 41370
rect 4408 41318 4418 41370
rect 4442 41318 4472 41370
rect 4472 41318 4498 41370
rect 4202 41316 4258 41318
rect 4282 41316 4338 41318
rect 4362 41316 4418 41318
rect 4442 41316 4498 41318
rect 4202 40282 4258 40284
rect 4282 40282 4338 40284
rect 4362 40282 4418 40284
rect 4442 40282 4498 40284
rect 4202 40230 4228 40282
rect 4228 40230 4258 40282
rect 4282 40230 4292 40282
rect 4292 40230 4338 40282
rect 4362 40230 4408 40282
rect 4408 40230 4418 40282
rect 4442 40230 4472 40282
rect 4472 40230 4498 40282
rect 4202 40228 4258 40230
rect 4282 40228 4338 40230
rect 4362 40228 4418 40230
rect 4442 40228 4498 40230
rect 4202 39194 4258 39196
rect 4282 39194 4338 39196
rect 4362 39194 4418 39196
rect 4442 39194 4498 39196
rect 4202 39142 4228 39194
rect 4228 39142 4258 39194
rect 4282 39142 4292 39194
rect 4292 39142 4338 39194
rect 4362 39142 4408 39194
rect 4408 39142 4418 39194
rect 4442 39142 4472 39194
rect 4472 39142 4498 39194
rect 4202 39140 4258 39142
rect 4282 39140 4338 39142
rect 4362 39140 4418 39142
rect 4442 39140 4498 39142
rect 4202 38106 4258 38108
rect 4282 38106 4338 38108
rect 4362 38106 4418 38108
rect 4442 38106 4498 38108
rect 4202 38054 4228 38106
rect 4228 38054 4258 38106
rect 4282 38054 4292 38106
rect 4292 38054 4338 38106
rect 4362 38054 4408 38106
rect 4408 38054 4418 38106
rect 4442 38054 4472 38106
rect 4472 38054 4498 38106
rect 4202 38052 4258 38054
rect 4282 38052 4338 38054
rect 4362 38052 4418 38054
rect 4442 38052 4498 38054
rect 4202 37018 4258 37020
rect 4282 37018 4338 37020
rect 4362 37018 4418 37020
rect 4442 37018 4498 37020
rect 4202 36966 4228 37018
rect 4228 36966 4258 37018
rect 4282 36966 4292 37018
rect 4292 36966 4338 37018
rect 4362 36966 4408 37018
rect 4408 36966 4418 37018
rect 4442 36966 4472 37018
rect 4472 36966 4498 37018
rect 4202 36964 4258 36966
rect 4282 36964 4338 36966
rect 4362 36964 4418 36966
rect 4442 36964 4498 36966
rect 4202 35930 4258 35932
rect 4282 35930 4338 35932
rect 4362 35930 4418 35932
rect 4442 35930 4498 35932
rect 4202 35878 4228 35930
rect 4228 35878 4258 35930
rect 4282 35878 4292 35930
rect 4292 35878 4338 35930
rect 4362 35878 4408 35930
rect 4408 35878 4418 35930
rect 4442 35878 4472 35930
rect 4472 35878 4498 35930
rect 4202 35876 4258 35878
rect 4282 35876 4338 35878
rect 4362 35876 4418 35878
rect 4442 35876 4498 35878
rect 4202 34842 4258 34844
rect 4282 34842 4338 34844
rect 4362 34842 4418 34844
rect 4442 34842 4498 34844
rect 4202 34790 4228 34842
rect 4228 34790 4258 34842
rect 4282 34790 4292 34842
rect 4292 34790 4338 34842
rect 4362 34790 4408 34842
rect 4408 34790 4418 34842
rect 4442 34790 4472 34842
rect 4472 34790 4498 34842
rect 4202 34788 4258 34790
rect 4282 34788 4338 34790
rect 4362 34788 4418 34790
rect 4442 34788 4498 34790
rect 4202 33754 4258 33756
rect 4282 33754 4338 33756
rect 4362 33754 4418 33756
rect 4442 33754 4498 33756
rect 4202 33702 4228 33754
rect 4228 33702 4258 33754
rect 4282 33702 4292 33754
rect 4292 33702 4338 33754
rect 4362 33702 4408 33754
rect 4408 33702 4418 33754
rect 4442 33702 4472 33754
rect 4472 33702 4498 33754
rect 4202 33700 4258 33702
rect 4282 33700 4338 33702
rect 4362 33700 4418 33702
rect 4442 33700 4498 33702
rect 4202 32666 4258 32668
rect 4282 32666 4338 32668
rect 4362 32666 4418 32668
rect 4442 32666 4498 32668
rect 4202 32614 4228 32666
rect 4228 32614 4258 32666
rect 4282 32614 4292 32666
rect 4292 32614 4338 32666
rect 4362 32614 4408 32666
rect 4408 32614 4418 32666
rect 4442 32614 4472 32666
rect 4472 32614 4498 32666
rect 4202 32612 4258 32614
rect 4282 32612 4338 32614
rect 4362 32612 4418 32614
rect 4442 32612 4498 32614
rect 4202 31578 4258 31580
rect 4282 31578 4338 31580
rect 4362 31578 4418 31580
rect 4442 31578 4498 31580
rect 4202 31526 4228 31578
rect 4228 31526 4258 31578
rect 4282 31526 4292 31578
rect 4292 31526 4338 31578
rect 4362 31526 4408 31578
rect 4408 31526 4418 31578
rect 4442 31526 4472 31578
rect 4472 31526 4498 31578
rect 4202 31524 4258 31526
rect 4282 31524 4338 31526
rect 4362 31524 4418 31526
rect 4442 31524 4498 31526
rect 4202 30490 4258 30492
rect 4282 30490 4338 30492
rect 4362 30490 4418 30492
rect 4442 30490 4498 30492
rect 4202 30438 4228 30490
rect 4228 30438 4258 30490
rect 4282 30438 4292 30490
rect 4292 30438 4338 30490
rect 4362 30438 4408 30490
rect 4408 30438 4418 30490
rect 4442 30438 4472 30490
rect 4472 30438 4498 30490
rect 4202 30436 4258 30438
rect 4282 30436 4338 30438
rect 4362 30436 4418 30438
rect 4442 30436 4498 30438
rect 4202 29402 4258 29404
rect 4282 29402 4338 29404
rect 4362 29402 4418 29404
rect 4442 29402 4498 29404
rect 4202 29350 4228 29402
rect 4228 29350 4258 29402
rect 4282 29350 4292 29402
rect 4292 29350 4338 29402
rect 4362 29350 4408 29402
rect 4408 29350 4418 29402
rect 4442 29350 4472 29402
rect 4472 29350 4498 29402
rect 4202 29348 4258 29350
rect 4282 29348 4338 29350
rect 4362 29348 4418 29350
rect 4442 29348 4498 29350
rect 4202 28314 4258 28316
rect 4282 28314 4338 28316
rect 4362 28314 4418 28316
rect 4442 28314 4498 28316
rect 4202 28262 4228 28314
rect 4228 28262 4258 28314
rect 4282 28262 4292 28314
rect 4292 28262 4338 28314
rect 4362 28262 4408 28314
rect 4408 28262 4418 28314
rect 4442 28262 4472 28314
rect 4472 28262 4498 28314
rect 4202 28260 4258 28262
rect 4282 28260 4338 28262
rect 4362 28260 4418 28262
rect 4442 28260 4498 28262
rect 4202 27226 4258 27228
rect 4282 27226 4338 27228
rect 4362 27226 4418 27228
rect 4442 27226 4498 27228
rect 4202 27174 4228 27226
rect 4228 27174 4258 27226
rect 4282 27174 4292 27226
rect 4292 27174 4338 27226
rect 4362 27174 4408 27226
rect 4408 27174 4418 27226
rect 4442 27174 4472 27226
rect 4472 27174 4498 27226
rect 4202 27172 4258 27174
rect 4282 27172 4338 27174
rect 4362 27172 4418 27174
rect 4442 27172 4498 27174
rect 4202 26138 4258 26140
rect 4282 26138 4338 26140
rect 4362 26138 4418 26140
rect 4442 26138 4498 26140
rect 4202 26086 4228 26138
rect 4228 26086 4258 26138
rect 4282 26086 4292 26138
rect 4292 26086 4338 26138
rect 4362 26086 4408 26138
rect 4408 26086 4418 26138
rect 4442 26086 4472 26138
rect 4472 26086 4498 26138
rect 4202 26084 4258 26086
rect 4282 26084 4338 26086
rect 4362 26084 4418 26086
rect 4442 26084 4498 26086
rect 4202 25050 4258 25052
rect 4282 25050 4338 25052
rect 4362 25050 4418 25052
rect 4442 25050 4498 25052
rect 4202 24998 4228 25050
rect 4228 24998 4258 25050
rect 4282 24998 4292 25050
rect 4292 24998 4338 25050
rect 4362 24998 4408 25050
rect 4408 24998 4418 25050
rect 4442 24998 4472 25050
rect 4472 24998 4498 25050
rect 4202 24996 4258 24998
rect 4282 24996 4338 24998
rect 4362 24996 4418 24998
rect 4442 24996 4498 24998
rect 4202 23962 4258 23964
rect 4282 23962 4338 23964
rect 4362 23962 4418 23964
rect 4442 23962 4498 23964
rect 4202 23910 4228 23962
rect 4228 23910 4258 23962
rect 4282 23910 4292 23962
rect 4292 23910 4338 23962
rect 4362 23910 4408 23962
rect 4408 23910 4418 23962
rect 4442 23910 4472 23962
rect 4472 23910 4498 23962
rect 4202 23908 4258 23910
rect 4282 23908 4338 23910
rect 4362 23908 4418 23910
rect 4442 23908 4498 23910
rect 4202 22874 4258 22876
rect 4282 22874 4338 22876
rect 4362 22874 4418 22876
rect 4442 22874 4498 22876
rect 4202 22822 4228 22874
rect 4228 22822 4258 22874
rect 4282 22822 4292 22874
rect 4292 22822 4338 22874
rect 4362 22822 4408 22874
rect 4408 22822 4418 22874
rect 4442 22822 4472 22874
rect 4472 22822 4498 22874
rect 4202 22820 4258 22822
rect 4282 22820 4338 22822
rect 4362 22820 4418 22822
rect 4442 22820 4498 22822
rect 4202 21786 4258 21788
rect 4282 21786 4338 21788
rect 4362 21786 4418 21788
rect 4442 21786 4498 21788
rect 4202 21734 4228 21786
rect 4228 21734 4258 21786
rect 4282 21734 4292 21786
rect 4292 21734 4338 21786
rect 4362 21734 4408 21786
rect 4408 21734 4418 21786
rect 4442 21734 4472 21786
rect 4472 21734 4498 21786
rect 4202 21732 4258 21734
rect 4282 21732 4338 21734
rect 4362 21732 4418 21734
rect 4442 21732 4498 21734
rect 4202 20698 4258 20700
rect 4282 20698 4338 20700
rect 4362 20698 4418 20700
rect 4442 20698 4498 20700
rect 4202 20646 4228 20698
rect 4228 20646 4258 20698
rect 4282 20646 4292 20698
rect 4292 20646 4338 20698
rect 4362 20646 4408 20698
rect 4408 20646 4418 20698
rect 4442 20646 4472 20698
rect 4472 20646 4498 20698
rect 4202 20644 4258 20646
rect 4282 20644 4338 20646
rect 4362 20644 4418 20646
rect 4442 20644 4498 20646
rect 4202 19610 4258 19612
rect 4282 19610 4338 19612
rect 4362 19610 4418 19612
rect 4442 19610 4498 19612
rect 4202 19558 4228 19610
rect 4228 19558 4258 19610
rect 4282 19558 4292 19610
rect 4292 19558 4338 19610
rect 4362 19558 4408 19610
rect 4408 19558 4418 19610
rect 4442 19558 4472 19610
rect 4472 19558 4498 19610
rect 4202 19556 4258 19558
rect 4282 19556 4338 19558
rect 4362 19556 4418 19558
rect 4442 19556 4498 19558
rect 4202 18522 4258 18524
rect 4282 18522 4338 18524
rect 4362 18522 4418 18524
rect 4442 18522 4498 18524
rect 4202 18470 4228 18522
rect 4228 18470 4258 18522
rect 4282 18470 4292 18522
rect 4292 18470 4338 18522
rect 4362 18470 4408 18522
rect 4408 18470 4418 18522
rect 4442 18470 4472 18522
rect 4472 18470 4498 18522
rect 4202 18468 4258 18470
rect 4282 18468 4338 18470
rect 4362 18468 4418 18470
rect 4442 18468 4498 18470
rect 4202 17434 4258 17436
rect 4282 17434 4338 17436
rect 4362 17434 4418 17436
rect 4442 17434 4498 17436
rect 4202 17382 4228 17434
rect 4228 17382 4258 17434
rect 4282 17382 4292 17434
rect 4292 17382 4338 17434
rect 4362 17382 4408 17434
rect 4408 17382 4418 17434
rect 4442 17382 4472 17434
rect 4472 17382 4498 17434
rect 4202 17380 4258 17382
rect 4282 17380 4338 17382
rect 4362 17380 4418 17382
rect 4442 17380 4498 17382
rect 4202 16346 4258 16348
rect 4282 16346 4338 16348
rect 4362 16346 4418 16348
rect 4442 16346 4498 16348
rect 4202 16294 4228 16346
rect 4228 16294 4258 16346
rect 4282 16294 4292 16346
rect 4292 16294 4338 16346
rect 4362 16294 4408 16346
rect 4408 16294 4418 16346
rect 4442 16294 4472 16346
rect 4472 16294 4498 16346
rect 4202 16292 4258 16294
rect 4282 16292 4338 16294
rect 4362 16292 4418 16294
rect 4442 16292 4498 16294
rect 4202 15258 4258 15260
rect 4282 15258 4338 15260
rect 4362 15258 4418 15260
rect 4442 15258 4498 15260
rect 4202 15206 4228 15258
rect 4228 15206 4258 15258
rect 4282 15206 4292 15258
rect 4292 15206 4338 15258
rect 4362 15206 4408 15258
rect 4408 15206 4418 15258
rect 4442 15206 4472 15258
rect 4472 15206 4498 15258
rect 4202 15204 4258 15206
rect 4282 15204 4338 15206
rect 4362 15204 4418 15206
rect 4442 15204 4498 15206
rect 4202 14170 4258 14172
rect 4282 14170 4338 14172
rect 4362 14170 4418 14172
rect 4442 14170 4498 14172
rect 4202 14118 4228 14170
rect 4228 14118 4258 14170
rect 4282 14118 4292 14170
rect 4292 14118 4338 14170
rect 4362 14118 4408 14170
rect 4408 14118 4418 14170
rect 4442 14118 4472 14170
rect 4472 14118 4498 14170
rect 4202 14116 4258 14118
rect 4282 14116 4338 14118
rect 4362 14116 4418 14118
rect 4442 14116 4498 14118
rect 4202 13082 4258 13084
rect 4282 13082 4338 13084
rect 4362 13082 4418 13084
rect 4442 13082 4498 13084
rect 4202 13030 4228 13082
rect 4228 13030 4258 13082
rect 4282 13030 4292 13082
rect 4292 13030 4338 13082
rect 4362 13030 4408 13082
rect 4408 13030 4418 13082
rect 4442 13030 4472 13082
rect 4472 13030 4498 13082
rect 4202 13028 4258 13030
rect 4282 13028 4338 13030
rect 4362 13028 4418 13030
rect 4442 13028 4498 13030
rect 4202 11994 4258 11996
rect 4282 11994 4338 11996
rect 4362 11994 4418 11996
rect 4442 11994 4498 11996
rect 4202 11942 4228 11994
rect 4228 11942 4258 11994
rect 4282 11942 4292 11994
rect 4292 11942 4338 11994
rect 4362 11942 4408 11994
rect 4408 11942 4418 11994
rect 4442 11942 4472 11994
rect 4472 11942 4498 11994
rect 4202 11940 4258 11942
rect 4282 11940 4338 11942
rect 4362 11940 4418 11942
rect 4442 11940 4498 11942
rect 4202 10906 4258 10908
rect 4282 10906 4338 10908
rect 4362 10906 4418 10908
rect 4442 10906 4498 10908
rect 4202 10854 4228 10906
rect 4228 10854 4258 10906
rect 4282 10854 4292 10906
rect 4292 10854 4338 10906
rect 4362 10854 4408 10906
rect 4408 10854 4418 10906
rect 4442 10854 4472 10906
rect 4472 10854 4498 10906
rect 4202 10852 4258 10854
rect 4282 10852 4338 10854
rect 4362 10852 4418 10854
rect 4442 10852 4498 10854
rect 4202 9818 4258 9820
rect 4282 9818 4338 9820
rect 4362 9818 4418 9820
rect 4442 9818 4498 9820
rect 4202 9766 4228 9818
rect 4228 9766 4258 9818
rect 4282 9766 4292 9818
rect 4292 9766 4338 9818
rect 4362 9766 4408 9818
rect 4408 9766 4418 9818
rect 4442 9766 4472 9818
rect 4472 9766 4498 9818
rect 4202 9764 4258 9766
rect 4282 9764 4338 9766
rect 4362 9764 4418 9766
rect 4442 9764 4498 9766
rect 4202 8730 4258 8732
rect 4282 8730 4338 8732
rect 4362 8730 4418 8732
rect 4442 8730 4498 8732
rect 4202 8678 4228 8730
rect 4228 8678 4258 8730
rect 4282 8678 4292 8730
rect 4292 8678 4338 8730
rect 4362 8678 4408 8730
rect 4408 8678 4418 8730
rect 4442 8678 4472 8730
rect 4472 8678 4498 8730
rect 4202 8676 4258 8678
rect 4282 8676 4338 8678
rect 4362 8676 4418 8678
rect 4442 8676 4498 8678
rect 4202 7642 4258 7644
rect 4282 7642 4338 7644
rect 4362 7642 4418 7644
rect 4442 7642 4498 7644
rect 4202 7590 4228 7642
rect 4228 7590 4258 7642
rect 4282 7590 4292 7642
rect 4292 7590 4338 7642
rect 4362 7590 4408 7642
rect 4408 7590 4418 7642
rect 4442 7590 4472 7642
rect 4472 7590 4498 7642
rect 4202 7588 4258 7590
rect 4282 7588 4338 7590
rect 4362 7588 4418 7590
rect 4442 7588 4498 7590
rect 4202 6554 4258 6556
rect 4282 6554 4338 6556
rect 4362 6554 4418 6556
rect 4442 6554 4498 6556
rect 4202 6502 4228 6554
rect 4228 6502 4258 6554
rect 4282 6502 4292 6554
rect 4292 6502 4338 6554
rect 4362 6502 4408 6554
rect 4408 6502 4418 6554
rect 4442 6502 4472 6554
rect 4472 6502 4498 6554
rect 4202 6500 4258 6502
rect 4282 6500 4338 6502
rect 4362 6500 4418 6502
rect 4442 6500 4498 6502
rect 4202 5466 4258 5468
rect 4282 5466 4338 5468
rect 4362 5466 4418 5468
rect 4442 5466 4498 5468
rect 4202 5414 4228 5466
rect 4228 5414 4258 5466
rect 4282 5414 4292 5466
rect 4292 5414 4338 5466
rect 4362 5414 4408 5466
rect 4408 5414 4418 5466
rect 4442 5414 4472 5466
rect 4472 5414 4498 5466
rect 4202 5412 4258 5414
rect 4282 5412 4338 5414
rect 4362 5412 4418 5414
rect 4442 5412 4498 5414
rect 4202 4378 4258 4380
rect 4282 4378 4338 4380
rect 4362 4378 4418 4380
rect 4442 4378 4498 4380
rect 4202 4326 4228 4378
rect 4228 4326 4258 4378
rect 4282 4326 4292 4378
rect 4292 4326 4338 4378
rect 4362 4326 4408 4378
rect 4408 4326 4418 4378
rect 4442 4326 4472 4378
rect 4472 4326 4498 4378
rect 4202 4324 4258 4326
rect 4282 4324 4338 4326
rect 4362 4324 4418 4326
rect 4442 4324 4498 4326
rect 4202 3290 4258 3292
rect 4282 3290 4338 3292
rect 4362 3290 4418 3292
rect 4442 3290 4498 3292
rect 4202 3238 4228 3290
rect 4228 3238 4258 3290
rect 4282 3238 4292 3290
rect 4292 3238 4338 3290
rect 4362 3238 4408 3290
rect 4408 3238 4418 3290
rect 4442 3238 4472 3290
rect 4472 3238 4498 3290
rect 4202 3236 4258 3238
rect 4282 3236 4338 3238
rect 4362 3236 4418 3238
rect 4442 3236 4498 3238
rect 4202 2202 4258 2204
rect 4282 2202 4338 2204
rect 4362 2202 4418 2204
rect 4442 2202 4498 2204
rect 4202 2150 4228 2202
rect 4228 2150 4258 2202
rect 4282 2150 4292 2202
rect 4292 2150 4338 2202
rect 4362 2150 4408 2202
rect 4408 2150 4418 2202
rect 4442 2150 4472 2202
rect 4472 2150 4498 2202
rect 4202 2148 4258 2150
rect 4282 2148 4338 2150
rect 4362 2148 4418 2150
rect 4442 2148 4498 2150
rect 5796 12008 5852 12064
rect 6808 12044 6810 12064
rect 6810 12044 6862 12064
rect 6862 12044 6864 12064
rect 6808 12008 6864 12044
rect 7728 3984 7784 4040
rect 8004 13812 8006 13832
rect 8006 13812 8058 13832
rect 8058 13812 8060 13832
rect 8004 13776 8060 13812
rect 8188 19116 8190 19136
rect 8190 19116 8242 19136
rect 8242 19116 8244 19136
rect 8188 19080 8244 19116
rect 8096 11756 8152 11792
rect 8096 11736 8098 11756
rect 8098 11736 8150 11756
rect 8150 11736 8152 11756
rect 8464 19352 8520 19408
rect 8924 19116 8926 19136
rect 8926 19116 8978 19136
rect 8978 19116 8980 19136
rect 8924 19080 8980 19116
rect 9200 17176 9256 17232
rect 9200 3032 9256 3088
rect 11132 3576 11188 3632
rect 11684 11736 11740 11792
rect 11224 3440 11280 3496
rect 12512 13812 12514 13832
rect 12514 13812 12566 13832
rect 12566 13812 12568 13832
rect 12512 13776 12568 13812
rect 14352 3712 14408 3768
rect 15180 15852 15182 15872
rect 15182 15852 15234 15872
rect 15234 15852 15236 15872
rect 15180 15816 15236 15852
rect 15180 11736 15236 11792
rect 15548 19352 15604 19408
rect 18492 55800 18548 55856
rect 18124 3304 18180 3360
rect 18216 3168 18272 3224
rect 19562 57146 19618 57148
rect 19642 57146 19698 57148
rect 19722 57146 19778 57148
rect 19802 57146 19858 57148
rect 19562 57094 19588 57146
rect 19588 57094 19618 57146
rect 19642 57094 19652 57146
rect 19652 57094 19698 57146
rect 19722 57094 19768 57146
rect 19768 57094 19778 57146
rect 19802 57094 19832 57146
rect 19832 57094 19858 57146
rect 19562 57092 19618 57094
rect 19642 57092 19698 57094
rect 19722 57092 19778 57094
rect 19802 57092 19858 57094
rect 19562 56058 19618 56060
rect 19642 56058 19698 56060
rect 19722 56058 19778 56060
rect 19802 56058 19858 56060
rect 19562 56006 19588 56058
rect 19588 56006 19618 56058
rect 19642 56006 19652 56058
rect 19652 56006 19698 56058
rect 19722 56006 19768 56058
rect 19768 56006 19778 56058
rect 19802 56006 19832 56058
rect 19832 56006 19858 56058
rect 19562 56004 19618 56006
rect 19642 56004 19698 56006
rect 19722 56004 19778 56006
rect 19802 56004 19858 56006
rect 19320 54596 19376 54632
rect 19320 54576 19322 54596
rect 19322 54576 19374 54596
rect 19374 54576 19376 54596
rect 18860 29008 18916 29064
rect 19562 54970 19618 54972
rect 19642 54970 19698 54972
rect 19722 54970 19778 54972
rect 19802 54970 19858 54972
rect 19562 54918 19588 54970
rect 19588 54918 19618 54970
rect 19642 54918 19652 54970
rect 19652 54918 19698 54970
rect 19722 54918 19768 54970
rect 19768 54918 19778 54970
rect 19802 54918 19832 54970
rect 19832 54918 19858 54970
rect 19562 54916 19618 54918
rect 19642 54916 19698 54918
rect 19722 54916 19778 54918
rect 19802 54916 19858 54918
rect 19562 53882 19618 53884
rect 19642 53882 19698 53884
rect 19722 53882 19778 53884
rect 19802 53882 19858 53884
rect 19562 53830 19588 53882
rect 19588 53830 19618 53882
rect 19642 53830 19652 53882
rect 19652 53830 19698 53882
rect 19722 53830 19768 53882
rect 19768 53830 19778 53882
rect 19802 53830 19832 53882
rect 19832 53830 19858 53882
rect 19562 53828 19618 53830
rect 19642 53828 19698 53830
rect 19722 53828 19778 53830
rect 19802 53828 19858 53830
rect 19562 52794 19618 52796
rect 19642 52794 19698 52796
rect 19722 52794 19778 52796
rect 19802 52794 19858 52796
rect 19562 52742 19588 52794
rect 19588 52742 19618 52794
rect 19642 52742 19652 52794
rect 19652 52742 19698 52794
rect 19722 52742 19768 52794
rect 19768 52742 19778 52794
rect 19802 52742 19832 52794
rect 19832 52742 19858 52794
rect 19562 52740 19618 52742
rect 19642 52740 19698 52742
rect 19722 52740 19778 52742
rect 19802 52740 19858 52742
rect 19562 51706 19618 51708
rect 19642 51706 19698 51708
rect 19722 51706 19778 51708
rect 19802 51706 19858 51708
rect 19562 51654 19588 51706
rect 19588 51654 19618 51706
rect 19642 51654 19652 51706
rect 19652 51654 19698 51706
rect 19722 51654 19768 51706
rect 19768 51654 19778 51706
rect 19802 51654 19832 51706
rect 19832 51654 19858 51706
rect 19562 51652 19618 51654
rect 19642 51652 19698 51654
rect 19722 51652 19778 51654
rect 19802 51652 19858 51654
rect 19562 50618 19618 50620
rect 19642 50618 19698 50620
rect 19722 50618 19778 50620
rect 19802 50618 19858 50620
rect 19562 50566 19588 50618
rect 19588 50566 19618 50618
rect 19642 50566 19652 50618
rect 19652 50566 19698 50618
rect 19722 50566 19768 50618
rect 19768 50566 19778 50618
rect 19802 50566 19832 50618
rect 19832 50566 19858 50618
rect 19562 50564 19618 50566
rect 19642 50564 19698 50566
rect 19722 50564 19778 50566
rect 19802 50564 19858 50566
rect 19562 49530 19618 49532
rect 19642 49530 19698 49532
rect 19722 49530 19778 49532
rect 19802 49530 19858 49532
rect 19562 49478 19588 49530
rect 19588 49478 19618 49530
rect 19642 49478 19652 49530
rect 19652 49478 19698 49530
rect 19722 49478 19768 49530
rect 19768 49478 19778 49530
rect 19802 49478 19832 49530
rect 19832 49478 19858 49530
rect 19562 49476 19618 49478
rect 19642 49476 19698 49478
rect 19722 49476 19778 49478
rect 19802 49476 19858 49478
rect 19562 48442 19618 48444
rect 19642 48442 19698 48444
rect 19722 48442 19778 48444
rect 19802 48442 19858 48444
rect 19562 48390 19588 48442
rect 19588 48390 19618 48442
rect 19642 48390 19652 48442
rect 19652 48390 19698 48442
rect 19722 48390 19768 48442
rect 19768 48390 19778 48442
rect 19802 48390 19832 48442
rect 19832 48390 19858 48442
rect 19562 48388 19618 48390
rect 19642 48388 19698 48390
rect 19722 48388 19778 48390
rect 19802 48388 19858 48390
rect 19562 47354 19618 47356
rect 19642 47354 19698 47356
rect 19722 47354 19778 47356
rect 19802 47354 19858 47356
rect 19562 47302 19588 47354
rect 19588 47302 19618 47354
rect 19642 47302 19652 47354
rect 19652 47302 19698 47354
rect 19722 47302 19768 47354
rect 19768 47302 19778 47354
rect 19802 47302 19832 47354
rect 19832 47302 19858 47354
rect 19562 47300 19618 47302
rect 19642 47300 19698 47302
rect 19722 47300 19778 47302
rect 19802 47300 19858 47302
rect 19562 46266 19618 46268
rect 19642 46266 19698 46268
rect 19722 46266 19778 46268
rect 19802 46266 19858 46268
rect 19562 46214 19588 46266
rect 19588 46214 19618 46266
rect 19642 46214 19652 46266
rect 19652 46214 19698 46266
rect 19722 46214 19768 46266
rect 19768 46214 19778 46266
rect 19802 46214 19832 46266
rect 19832 46214 19858 46266
rect 19562 46212 19618 46214
rect 19642 46212 19698 46214
rect 19722 46212 19778 46214
rect 19802 46212 19858 46214
rect 19562 45178 19618 45180
rect 19642 45178 19698 45180
rect 19722 45178 19778 45180
rect 19802 45178 19858 45180
rect 19562 45126 19588 45178
rect 19588 45126 19618 45178
rect 19642 45126 19652 45178
rect 19652 45126 19698 45178
rect 19722 45126 19768 45178
rect 19768 45126 19778 45178
rect 19802 45126 19832 45178
rect 19832 45126 19858 45178
rect 19562 45124 19618 45126
rect 19642 45124 19698 45126
rect 19722 45124 19778 45126
rect 19802 45124 19858 45126
rect 19562 44090 19618 44092
rect 19642 44090 19698 44092
rect 19722 44090 19778 44092
rect 19802 44090 19858 44092
rect 19562 44038 19588 44090
rect 19588 44038 19618 44090
rect 19642 44038 19652 44090
rect 19652 44038 19698 44090
rect 19722 44038 19768 44090
rect 19768 44038 19778 44090
rect 19802 44038 19832 44090
rect 19832 44038 19858 44090
rect 19562 44036 19618 44038
rect 19642 44036 19698 44038
rect 19722 44036 19778 44038
rect 19802 44036 19858 44038
rect 19562 43002 19618 43004
rect 19642 43002 19698 43004
rect 19722 43002 19778 43004
rect 19802 43002 19858 43004
rect 19562 42950 19588 43002
rect 19588 42950 19618 43002
rect 19642 42950 19652 43002
rect 19652 42950 19698 43002
rect 19722 42950 19768 43002
rect 19768 42950 19778 43002
rect 19802 42950 19832 43002
rect 19832 42950 19858 43002
rect 19562 42948 19618 42950
rect 19642 42948 19698 42950
rect 19722 42948 19778 42950
rect 19802 42948 19858 42950
rect 19562 41914 19618 41916
rect 19642 41914 19698 41916
rect 19722 41914 19778 41916
rect 19802 41914 19858 41916
rect 19562 41862 19588 41914
rect 19588 41862 19618 41914
rect 19642 41862 19652 41914
rect 19652 41862 19698 41914
rect 19722 41862 19768 41914
rect 19768 41862 19778 41914
rect 19802 41862 19832 41914
rect 19832 41862 19858 41914
rect 19562 41860 19618 41862
rect 19642 41860 19698 41862
rect 19722 41860 19778 41862
rect 19802 41860 19858 41862
rect 19562 40826 19618 40828
rect 19642 40826 19698 40828
rect 19722 40826 19778 40828
rect 19802 40826 19858 40828
rect 19562 40774 19588 40826
rect 19588 40774 19618 40826
rect 19642 40774 19652 40826
rect 19652 40774 19698 40826
rect 19722 40774 19768 40826
rect 19768 40774 19778 40826
rect 19802 40774 19832 40826
rect 19832 40774 19858 40826
rect 19562 40772 19618 40774
rect 19642 40772 19698 40774
rect 19722 40772 19778 40774
rect 19802 40772 19858 40774
rect 19562 39738 19618 39740
rect 19642 39738 19698 39740
rect 19722 39738 19778 39740
rect 19802 39738 19858 39740
rect 19562 39686 19588 39738
rect 19588 39686 19618 39738
rect 19642 39686 19652 39738
rect 19652 39686 19698 39738
rect 19722 39686 19768 39738
rect 19768 39686 19778 39738
rect 19802 39686 19832 39738
rect 19832 39686 19858 39738
rect 19562 39684 19618 39686
rect 19642 39684 19698 39686
rect 19722 39684 19778 39686
rect 19802 39684 19858 39686
rect 19562 38650 19618 38652
rect 19642 38650 19698 38652
rect 19722 38650 19778 38652
rect 19802 38650 19858 38652
rect 19562 38598 19588 38650
rect 19588 38598 19618 38650
rect 19642 38598 19652 38650
rect 19652 38598 19698 38650
rect 19722 38598 19768 38650
rect 19768 38598 19778 38650
rect 19802 38598 19832 38650
rect 19832 38598 19858 38650
rect 19562 38596 19618 38598
rect 19642 38596 19698 38598
rect 19722 38596 19778 38598
rect 19802 38596 19858 38598
rect 19562 37562 19618 37564
rect 19642 37562 19698 37564
rect 19722 37562 19778 37564
rect 19802 37562 19858 37564
rect 19562 37510 19588 37562
rect 19588 37510 19618 37562
rect 19642 37510 19652 37562
rect 19652 37510 19698 37562
rect 19722 37510 19768 37562
rect 19768 37510 19778 37562
rect 19802 37510 19832 37562
rect 19832 37510 19858 37562
rect 19562 37508 19618 37510
rect 19642 37508 19698 37510
rect 19722 37508 19778 37510
rect 19802 37508 19858 37510
rect 19562 36474 19618 36476
rect 19642 36474 19698 36476
rect 19722 36474 19778 36476
rect 19802 36474 19858 36476
rect 19562 36422 19588 36474
rect 19588 36422 19618 36474
rect 19642 36422 19652 36474
rect 19652 36422 19698 36474
rect 19722 36422 19768 36474
rect 19768 36422 19778 36474
rect 19802 36422 19832 36474
rect 19832 36422 19858 36474
rect 19562 36420 19618 36422
rect 19642 36420 19698 36422
rect 19722 36420 19778 36422
rect 19802 36420 19858 36422
rect 19562 35386 19618 35388
rect 19642 35386 19698 35388
rect 19722 35386 19778 35388
rect 19802 35386 19858 35388
rect 19562 35334 19588 35386
rect 19588 35334 19618 35386
rect 19642 35334 19652 35386
rect 19652 35334 19698 35386
rect 19722 35334 19768 35386
rect 19768 35334 19778 35386
rect 19802 35334 19832 35386
rect 19832 35334 19858 35386
rect 19562 35332 19618 35334
rect 19642 35332 19698 35334
rect 19722 35332 19778 35334
rect 19802 35332 19858 35334
rect 19562 34298 19618 34300
rect 19642 34298 19698 34300
rect 19722 34298 19778 34300
rect 19802 34298 19858 34300
rect 19562 34246 19588 34298
rect 19588 34246 19618 34298
rect 19642 34246 19652 34298
rect 19652 34246 19698 34298
rect 19722 34246 19768 34298
rect 19768 34246 19778 34298
rect 19802 34246 19832 34298
rect 19832 34246 19858 34298
rect 19562 34244 19618 34246
rect 19642 34244 19698 34246
rect 19722 34244 19778 34246
rect 19802 34244 19858 34246
rect 19562 33210 19618 33212
rect 19642 33210 19698 33212
rect 19722 33210 19778 33212
rect 19802 33210 19858 33212
rect 19562 33158 19588 33210
rect 19588 33158 19618 33210
rect 19642 33158 19652 33210
rect 19652 33158 19698 33210
rect 19722 33158 19768 33210
rect 19768 33158 19778 33210
rect 19802 33158 19832 33210
rect 19832 33158 19858 33210
rect 19562 33156 19618 33158
rect 19642 33156 19698 33158
rect 19722 33156 19778 33158
rect 19802 33156 19858 33158
rect 19562 32122 19618 32124
rect 19642 32122 19698 32124
rect 19722 32122 19778 32124
rect 19802 32122 19858 32124
rect 19562 32070 19588 32122
rect 19588 32070 19618 32122
rect 19642 32070 19652 32122
rect 19652 32070 19698 32122
rect 19722 32070 19768 32122
rect 19768 32070 19778 32122
rect 19802 32070 19832 32122
rect 19832 32070 19858 32122
rect 19562 32068 19618 32070
rect 19642 32068 19698 32070
rect 19722 32068 19778 32070
rect 19802 32068 19858 32070
rect 19562 31034 19618 31036
rect 19642 31034 19698 31036
rect 19722 31034 19778 31036
rect 19802 31034 19858 31036
rect 19562 30982 19588 31034
rect 19588 30982 19618 31034
rect 19642 30982 19652 31034
rect 19652 30982 19698 31034
rect 19722 30982 19768 31034
rect 19768 30982 19778 31034
rect 19802 30982 19832 31034
rect 19832 30982 19858 31034
rect 19562 30980 19618 30982
rect 19642 30980 19698 30982
rect 19722 30980 19778 30982
rect 19802 30980 19858 30982
rect 19562 29946 19618 29948
rect 19642 29946 19698 29948
rect 19722 29946 19778 29948
rect 19802 29946 19858 29948
rect 19562 29894 19588 29946
rect 19588 29894 19618 29946
rect 19642 29894 19652 29946
rect 19652 29894 19698 29946
rect 19722 29894 19768 29946
rect 19768 29894 19778 29946
rect 19802 29894 19832 29946
rect 19832 29894 19858 29946
rect 19562 29892 19618 29894
rect 19642 29892 19698 29894
rect 19722 29892 19778 29894
rect 19802 29892 19858 29894
rect 18952 28872 19008 28928
rect 19562 28858 19618 28860
rect 19642 28858 19698 28860
rect 19722 28858 19778 28860
rect 19802 28858 19858 28860
rect 19562 28806 19588 28858
rect 19588 28806 19618 28858
rect 19642 28806 19652 28858
rect 19652 28806 19698 28858
rect 19722 28806 19768 28858
rect 19768 28806 19778 28858
rect 19802 28806 19832 28858
rect 19832 28806 19858 28858
rect 19562 28804 19618 28806
rect 19642 28804 19698 28806
rect 19722 28804 19778 28806
rect 19802 28804 19858 28806
rect 19562 27770 19618 27772
rect 19642 27770 19698 27772
rect 19722 27770 19778 27772
rect 19802 27770 19858 27772
rect 19562 27718 19588 27770
rect 19588 27718 19618 27770
rect 19642 27718 19652 27770
rect 19652 27718 19698 27770
rect 19722 27718 19768 27770
rect 19768 27718 19778 27770
rect 19802 27718 19832 27770
rect 19832 27718 19858 27770
rect 19562 27716 19618 27718
rect 19642 27716 19698 27718
rect 19722 27716 19778 27718
rect 19802 27716 19858 27718
rect 19562 26682 19618 26684
rect 19642 26682 19698 26684
rect 19722 26682 19778 26684
rect 19802 26682 19858 26684
rect 19562 26630 19588 26682
rect 19588 26630 19618 26682
rect 19642 26630 19652 26682
rect 19652 26630 19698 26682
rect 19722 26630 19768 26682
rect 19768 26630 19778 26682
rect 19802 26630 19832 26682
rect 19832 26630 19858 26682
rect 19562 26628 19618 26630
rect 19642 26628 19698 26630
rect 19722 26628 19778 26630
rect 19802 26628 19858 26630
rect 19562 25594 19618 25596
rect 19642 25594 19698 25596
rect 19722 25594 19778 25596
rect 19802 25594 19858 25596
rect 19562 25542 19588 25594
rect 19588 25542 19618 25594
rect 19642 25542 19652 25594
rect 19652 25542 19698 25594
rect 19722 25542 19768 25594
rect 19768 25542 19778 25594
rect 19802 25542 19832 25594
rect 19832 25542 19858 25594
rect 19562 25540 19618 25542
rect 19642 25540 19698 25542
rect 19722 25540 19778 25542
rect 19802 25540 19858 25542
rect 19562 24506 19618 24508
rect 19642 24506 19698 24508
rect 19722 24506 19778 24508
rect 19802 24506 19858 24508
rect 19562 24454 19588 24506
rect 19588 24454 19618 24506
rect 19642 24454 19652 24506
rect 19652 24454 19698 24506
rect 19722 24454 19768 24506
rect 19768 24454 19778 24506
rect 19802 24454 19832 24506
rect 19832 24454 19858 24506
rect 19562 24452 19618 24454
rect 19642 24452 19698 24454
rect 19722 24452 19778 24454
rect 19802 24452 19858 24454
rect 18860 17992 18916 18048
rect 18952 17856 19008 17912
rect 18952 3712 19008 3768
rect 19562 23418 19618 23420
rect 19642 23418 19698 23420
rect 19722 23418 19778 23420
rect 19802 23418 19858 23420
rect 19562 23366 19588 23418
rect 19588 23366 19618 23418
rect 19642 23366 19652 23418
rect 19652 23366 19698 23418
rect 19722 23366 19768 23418
rect 19768 23366 19778 23418
rect 19802 23366 19832 23418
rect 19832 23366 19858 23418
rect 19562 23364 19618 23366
rect 19642 23364 19698 23366
rect 19722 23364 19778 23366
rect 19802 23364 19858 23366
rect 19562 22330 19618 22332
rect 19642 22330 19698 22332
rect 19722 22330 19778 22332
rect 19802 22330 19858 22332
rect 19562 22278 19588 22330
rect 19588 22278 19618 22330
rect 19642 22278 19652 22330
rect 19652 22278 19698 22330
rect 19722 22278 19768 22330
rect 19768 22278 19778 22330
rect 19802 22278 19832 22330
rect 19832 22278 19858 22330
rect 19562 22276 19618 22278
rect 19642 22276 19698 22278
rect 19722 22276 19778 22278
rect 19802 22276 19858 22278
rect 19562 21242 19618 21244
rect 19642 21242 19698 21244
rect 19722 21242 19778 21244
rect 19802 21242 19858 21244
rect 19562 21190 19588 21242
rect 19588 21190 19618 21242
rect 19642 21190 19652 21242
rect 19652 21190 19698 21242
rect 19722 21190 19768 21242
rect 19768 21190 19778 21242
rect 19802 21190 19832 21242
rect 19832 21190 19858 21242
rect 19562 21188 19618 21190
rect 19642 21188 19698 21190
rect 19722 21188 19778 21190
rect 19802 21188 19858 21190
rect 19562 20154 19618 20156
rect 19642 20154 19698 20156
rect 19722 20154 19778 20156
rect 19802 20154 19858 20156
rect 19562 20102 19588 20154
rect 19588 20102 19618 20154
rect 19642 20102 19652 20154
rect 19652 20102 19698 20154
rect 19722 20102 19768 20154
rect 19768 20102 19778 20154
rect 19802 20102 19832 20154
rect 19832 20102 19858 20154
rect 19562 20100 19618 20102
rect 19642 20100 19698 20102
rect 19722 20100 19778 20102
rect 19802 20100 19858 20102
rect 19562 19066 19618 19068
rect 19642 19066 19698 19068
rect 19722 19066 19778 19068
rect 19802 19066 19858 19068
rect 19562 19014 19588 19066
rect 19588 19014 19618 19066
rect 19642 19014 19652 19066
rect 19652 19014 19698 19066
rect 19722 19014 19768 19066
rect 19768 19014 19778 19066
rect 19802 19014 19832 19066
rect 19832 19014 19858 19066
rect 19562 19012 19618 19014
rect 19642 19012 19698 19014
rect 19722 19012 19778 19014
rect 19802 19012 19858 19014
rect 19562 17978 19618 17980
rect 19642 17978 19698 17980
rect 19722 17978 19778 17980
rect 19802 17978 19858 17980
rect 19562 17926 19588 17978
rect 19588 17926 19618 17978
rect 19642 17926 19652 17978
rect 19652 17926 19698 17978
rect 19722 17926 19768 17978
rect 19768 17926 19778 17978
rect 19802 17926 19832 17978
rect 19832 17926 19858 17978
rect 19562 17924 19618 17926
rect 19642 17924 19698 17926
rect 19722 17924 19778 17926
rect 19802 17924 19858 17926
rect 19320 17484 19322 17504
rect 19322 17484 19374 17504
rect 19374 17484 19376 17504
rect 19320 17448 19376 17484
rect 19562 16890 19618 16892
rect 19642 16890 19698 16892
rect 19722 16890 19778 16892
rect 19802 16890 19858 16892
rect 19562 16838 19588 16890
rect 19588 16838 19618 16890
rect 19642 16838 19652 16890
rect 19652 16838 19698 16890
rect 19722 16838 19768 16890
rect 19768 16838 19778 16890
rect 19802 16838 19832 16890
rect 19832 16838 19858 16890
rect 19562 16836 19618 16838
rect 19642 16836 19698 16838
rect 19722 16836 19778 16838
rect 19802 16836 19858 16838
rect 19562 15802 19618 15804
rect 19642 15802 19698 15804
rect 19722 15802 19778 15804
rect 19802 15802 19858 15804
rect 19562 15750 19588 15802
rect 19588 15750 19618 15802
rect 19642 15750 19652 15802
rect 19652 15750 19698 15802
rect 19722 15750 19768 15802
rect 19768 15750 19778 15802
rect 19802 15750 19832 15802
rect 19832 15750 19858 15802
rect 19562 15748 19618 15750
rect 19642 15748 19698 15750
rect 19722 15748 19778 15750
rect 19802 15748 19858 15750
rect 19562 14714 19618 14716
rect 19642 14714 19698 14716
rect 19722 14714 19778 14716
rect 19802 14714 19858 14716
rect 19562 14662 19588 14714
rect 19588 14662 19618 14714
rect 19642 14662 19652 14714
rect 19652 14662 19698 14714
rect 19722 14662 19768 14714
rect 19768 14662 19778 14714
rect 19802 14662 19832 14714
rect 19832 14662 19858 14714
rect 19562 14660 19618 14662
rect 19642 14660 19698 14662
rect 19722 14660 19778 14662
rect 19802 14660 19858 14662
rect 19562 13626 19618 13628
rect 19642 13626 19698 13628
rect 19722 13626 19778 13628
rect 19802 13626 19858 13628
rect 19562 13574 19588 13626
rect 19588 13574 19618 13626
rect 19642 13574 19652 13626
rect 19652 13574 19698 13626
rect 19722 13574 19768 13626
rect 19768 13574 19778 13626
rect 19802 13574 19832 13626
rect 19832 13574 19858 13626
rect 19562 13572 19618 13574
rect 19642 13572 19698 13574
rect 19722 13572 19778 13574
rect 19802 13572 19858 13574
rect 19562 12538 19618 12540
rect 19642 12538 19698 12540
rect 19722 12538 19778 12540
rect 19802 12538 19858 12540
rect 19562 12486 19588 12538
rect 19588 12486 19618 12538
rect 19642 12486 19652 12538
rect 19652 12486 19698 12538
rect 19722 12486 19768 12538
rect 19768 12486 19778 12538
rect 19802 12486 19832 12538
rect 19832 12486 19858 12538
rect 19562 12484 19618 12486
rect 19642 12484 19698 12486
rect 19722 12484 19778 12486
rect 19802 12484 19858 12486
rect 19562 11450 19618 11452
rect 19642 11450 19698 11452
rect 19722 11450 19778 11452
rect 19802 11450 19858 11452
rect 19562 11398 19588 11450
rect 19588 11398 19618 11450
rect 19642 11398 19652 11450
rect 19652 11398 19698 11450
rect 19722 11398 19768 11450
rect 19768 11398 19778 11450
rect 19802 11398 19832 11450
rect 19832 11398 19858 11450
rect 19562 11396 19618 11398
rect 19642 11396 19698 11398
rect 19722 11396 19778 11398
rect 19802 11396 19858 11398
rect 19562 10362 19618 10364
rect 19642 10362 19698 10364
rect 19722 10362 19778 10364
rect 19802 10362 19858 10364
rect 19562 10310 19588 10362
rect 19588 10310 19618 10362
rect 19642 10310 19652 10362
rect 19652 10310 19698 10362
rect 19722 10310 19768 10362
rect 19768 10310 19778 10362
rect 19802 10310 19832 10362
rect 19832 10310 19858 10362
rect 19562 10308 19618 10310
rect 19642 10308 19698 10310
rect 19722 10308 19778 10310
rect 19802 10308 19858 10310
rect 19562 9274 19618 9276
rect 19642 9274 19698 9276
rect 19722 9274 19778 9276
rect 19802 9274 19858 9276
rect 19562 9222 19588 9274
rect 19588 9222 19618 9274
rect 19642 9222 19652 9274
rect 19652 9222 19698 9274
rect 19722 9222 19768 9274
rect 19768 9222 19778 9274
rect 19802 9222 19832 9274
rect 19832 9222 19858 9274
rect 19562 9220 19618 9222
rect 19642 9220 19698 9222
rect 19722 9220 19778 9222
rect 19802 9220 19858 9222
rect 19562 8186 19618 8188
rect 19642 8186 19698 8188
rect 19722 8186 19778 8188
rect 19802 8186 19858 8188
rect 19562 8134 19588 8186
rect 19588 8134 19618 8186
rect 19642 8134 19652 8186
rect 19652 8134 19698 8186
rect 19722 8134 19768 8186
rect 19768 8134 19778 8186
rect 19802 8134 19832 8186
rect 19832 8134 19858 8186
rect 19562 8132 19618 8134
rect 19642 8132 19698 8134
rect 19722 8132 19778 8134
rect 19802 8132 19858 8134
rect 19872 7656 19928 7712
rect 19872 7520 19928 7576
rect 19562 7098 19618 7100
rect 19642 7098 19698 7100
rect 19722 7098 19778 7100
rect 19802 7098 19858 7100
rect 19562 7046 19588 7098
rect 19588 7046 19618 7098
rect 19642 7046 19652 7098
rect 19652 7046 19698 7098
rect 19722 7046 19768 7098
rect 19768 7046 19778 7098
rect 19802 7046 19832 7098
rect 19832 7046 19858 7098
rect 19562 7044 19618 7046
rect 19642 7044 19698 7046
rect 19722 7044 19778 7046
rect 19802 7044 19858 7046
rect 19562 6010 19618 6012
rect 19642 6010 19698 6012
rect 19722 6010 19778 6012
rect 19802 6010 19858 6012
rect 19562 5958 19588 6010
rect 19588 5958 19618 6010
rect 19642 5958 19652 6010
rect 19652 5958 19698 6010
rect 19722 5958 19768 6010
rect 19768 5958 19778 6010
rect 19802 5958 19832 6010
rect 19832 5958 19858 6010
rect 19562 5956 19618 5958
rect 19642 5956 19698 5958
rect 19722 5956 19778 5958
rect 19802 5956 19858 5958
rect 19562 4922 19618 4924
rect 19642 4922 19698 4924
rect 19722 4922 19778 4924
rect 19802 4922 19858 4924
rect 19562 4870 19588 4922
rect 19588 4870 19618 4922
rect 19642 4870 19652 4922
rect 19652 4870 19698 4922
rect 19722 4870 19768 4922
rect 19768 4870 19778 4922
rect 19802 4870 19832 4922
rect 19832 4870 19858 4922
rect 19562 4868 19618 4870
rect 19642 4868 19698 4870
rect 19722 4868 19778 4870
rect 19802 4868 19858 4870
rect 19562 3834 19618 3836
rect 19642 3834 19698 3836
rect 19722 3834 19778 3836
rect 19802 3834 19858 3836
rect 19562 3782 19588 3834
rect 19588 3782 19618 3834
rect 19642 3782 19652 3834
rect 19652 3782 19698 3834
rect 19722 3782 19768 3834
rect 19768 3782 19778 3834
rect 19802 3782 19832 3834
rect 19832 3782 19858 3834
rect 19562 3780 19618 3782
rect 19642 3780 19698 3782
rect 19722 3780 19778 3782
rect 19802 3780 19858 3782
rect 19562 2746 19618 2748
rect 19642 2746 19698 2748
rect 19722 2746 19778 2748
rect 19802 2746 19858 2748
rect 19562 2694 19588 2746
rect 19588 2694 19618 2746
rect 19642 2694 19652 2746
rect 19652 2694 19698 2746
rect 19722 2694 19768 2746
rect 19768 2694 19778 2746
rect 19802 2694 19832 2746
rect 19832 2694 19858 2746
rect 19562 2692 19618 2694
rect 19642 2692 19698 2694
rect 19722 2692 19778 2694
rect 19802 2692 19858 2694
rect 20148 7520 20204 7576
rect 20424 856 20480 912
rect 23000 44104 23056 44160
rect 23184 44104 23240 44160
rect 23552 54576 23608 54632
rect 24104 38664 24160 38720
rect 24104 38528 24160 38584
rect 23368 17176 23424 17232
rect 23276 15136 23332 15192
rect 23552 23296 23608 23352
rect 24564 17484 24566 17504
rect 24566 17484 24618 17504
rect 24618 17484 24620 17504
rect 24564 17448 24620 17484
rect 24748 15816 24804 15872
rect 24748 11600 24804 11656
rect 26956 56752 27012 56808
rect 26864 56616 26920 56672
rect 26680 56364 26736 56400
rect 26680 56344 26682 56364
rect 26682 56344 26734 56364
rect 26734 56344 26736 56364
rect 28152 56380 28154 56400
rect 28154 56380 28206 56400
rect 28206 56380 28208 56400
rect 28152 56344 28208 56380
rect 27416 55564 27418 55584
rect 27418 55564 27470 55584
rect 27470 55564 27472 55584
rect 27416 55528 27472 55564
rect 26864 3304 26920 3360
rect 26864 2760 26920 2816
rect 29348 38664 29404 38720
rect 29256 38528 29312 38584
rect 31188 55564 31190 55584
rect 31190 55564 31242 55584
rect 31242 55564 31244 55584
rect 31188 55528 31244 55564
rect 31648 56072 31704 56128
rect 31832 56072 31888 56128
rect 31556 55664 31612 55720
rect 31740 55664 31796 55720
rect 32476 56208 32532 56264
rect 31740 3884 31742 3904
rect 31742 3884 31794 3904
rect 31794 3884 31796 3904
rect 31740 3848 31796 3884
rect 31832 3304 31888 3360
rect 32476 3712 32532 3768
rect 33764 56344 33820 56400
rect 33028 3848 33084 3904
rect 33672 3304 33728 3360
rect 34922 57690 34978 57692
rect 35002 57690 35058 57692
rect 35082 57690 35138 57692
rect 35162 57690 35218 57692
rect 34922 57638 34948 57690
rect 34948 57638 34978 57690
rect 35002 57638 35012 57690
rect 35012 57638 35058 57690
rect 35082 57638 35128 57690
rect 35128 57638 35138 57690
rect 35162 57638 35192 57690
rect 35192 57638 35218 57690
rect 34922 57636 34978 57638
rect 35002 57636 35058 57638
rect 35082 57636 35138 57638
rect 35162 57636 35218 57638
rect 34922 56602 34978 56604
rect 35002 56602 35058 56604
rect 35082 56602 35138 56604
rect 35162 56602 35218 56604
rect 34922 56550 34948 56602
rect 34948 56550 34978 56602
rect 35002 56550 35012 56602
rect 35012 56550 35058 56602
rect 35082 56550 35128 56602
rect 35128 56550 35138 56602
rect 35162 56550 35192 56602
rect 35192 56550 35218 56602
rect 34922 56548 34978 56550
rect 35002 56548 35058 56550
rect 35082 56548 35138 56550
rect 35162 56548 35218 56550
rect 34922 55514 34978 55516
rect 35002 55514 35058 55516
rect 35082 55514 35138 55516
rect 35162 55514 35218 55516
rect 34922 55462 34948 55514
rect 34948 55462 34978 55514
rect 35002 55462 35012 55514
rect 35012 55462 35058 55514
rect 35082 55462 35128 55514
rect 35128 55462 35138 55514
rect 35162 55462 35192 55514
rect 35192 55462 35218 55514
rect 34922 55460 34978 55462
rect 35002 55460 35058 55462
rect 35082 55460 35138 55462
rect 35162 55460 35218 55462
rect 34922 54426 34978 54428
rect 35002 54426 35058 54428
rect 35082 54426 35138 54428
rect 35162 54426 35218 54428
rect 34922 54374 34948 54426
rect 34948 54374 34978 54426
rect 35002 54374 35012 54426
rect 35012 54374 35058 54426
rect 35082 54374 35128 54426
rect 35128 54374 35138 54426
rect 35162 54374 35192 54426
rect 35192 54374 35218 54426
rect 34922 54372 34978 54374
rect 35002 54372 35058 54374
rect 35082 54372 35138 54374
rect 35162 54372 35218 54374
rect 34922 53338 34978 53340
rect 35002 53338 35058 53340
rect 35082 53338 35138 53340
rect 35162 53338 35218 53340
rect 34922 53286 34948 53338
rect 34948 53286 34978 53338
rect 35002 53286 35012 53338
rect 35012 53286 35058 53338
rect 35082 53286 35128 53338
rect 35128 53286 35138 53338
rect 35162 53286 35192 53338
rect 35192 53286 35218 53338
rect 34922 53284 34978 53286
rect 35002 53284 35058 53286
rect 35082 53284 35138 53286
rect 35162 53284 35218 53286
rect 34922 52250 34978 52252
rect 35002 52250 35058 52252
rect 35082 52250 35138 52252
rect 35162 52250 35218 52252
rect 34922 52198 34948 52250
rect 34948 52198 34978 52250
rect 35002 52198 35012 52250
rect 35012 52198 35058 52250
rect 35082 52198 35128 52250
rect 35128 52198 35138 52250
rect 35162 52198 35192 52250
rect 35192 52198 35218 52250
rect 34922 52196 34978 52198
rect 35002 52196 35058 52198
rect 35082 52196 35138 52198
rect 35162 52196 35218 52198
rect 34922 51162 34978 51164
rect 35002 51162 35058 51164
rect 35082 51162 35138 51164
rect 35162 51162 35218 51164
rect 34922 51110 34948 51162
rect 34948 51110 34978 51162
rect 35002 51110 35012 51162
rect 35012 51110 35058 51162
rect 35082 51110 35128 51162
rect 35128 51110 35138 51162
rect 35162 51110 35192 51162
rect 35192 51110 35218 51162
rect 34922 51108 34978 51110
rect 35002 51108 35058 51110
rect 35082 51108 35138 51110
rect 35162 51108 35218 51110
rect 34922 50074 34978 50076
rect 35002 50074 35058 50076
rect 35082 50074 35138 50076
rect 35162 50074 35218 50076
rect 34922 50022 34948 50074
rect 34948 50022 34978 50074
rect 35002 50022 35012 50074
rect 35012 50022 35058 50074
rect 35082 50022 35128 50074
rect 35128 50022 35138 50074
rect 35162 50022 35192 50074
rect 35192 50022 35218 50074
rect 34922 50020 34978 50022
rect 35002 50020 35058 50022
rect 35082 50020 35138 50022
rect 35162 50020 35218 50022
rect 34922 48986 34978 48988
rect 35002 48986 35058 48988
rect 35082 48986 35138 48988
rect 35162 48986 35218 48988
rect 34922 48934 34948 48986
rect 34948 48934 34978 48986
rect 35002 48934 35012 48986
rect 35012 48934 35058 48986
rect 35082 48934 35128 48986
rect 35128 48934 35138 48986
rect 35162 48934 35192 48986
rect 35192 48934 35218 48986
rect 34922 48932 34978 48934
rect 35002 48932 35058 48934
rect 35082 48932 35138 48934
rect 35162 48932 35218 48934
rect 34922 47898 34978 47900
rect 35002 47898 35058 47900
rect 35082 47898 35138 47900
rect 35162 47898 35218 47900
rect 34922 47846 34948 47898
rect 34948 47846 34978 47898
rect 35002 47846 35012 47898
rect 35012 47846 35058 47898
rect 35082 47846 35128 47898
rect 35128 47846 35138 47898
rect 35162 47846 35192 47898
rect 35192 47846 35218 47898
rect 34922 47844 34978 47846
rect 35002 47844 35058 47846
rect 35082 47844 35138 47846
rect 35162 47844 35218 47846
rect 34922 46810 34978 46812
rect 35002 46810 35058 46812
rect 35082 46810 35138 46812
rect 35162 46810 35218 46812
rect 34922 46758 34948 46810
rect 34948 46758 34978 46810
rect 35002 46758 35012 46810
rect 35012 46758 35058 46810
rect 35082 46758 35128 46810
rect 35128 46758 35138 46810
rect 35162 46758 35192 46810
rect 35192 46758 35218 46810
rect 34922 46756 34978 46758
rect 35002 46756 35058 46758
rect 35082 46756 35138 46758
rect 35162 46756 35218 46758
rect 34922 45722 34978 45724
rect 35002 45722 35058 45724
rect 35082 45722 35138 45724
rect 35162 45722 35218 45724
rect 34922 45670 34948 45722
rect 34948 45670 34978 45722
rect 35002 45670 35012 45722
rect 35012 45670 35058 45722
rect 35082 45670 35128 45722
rect 35128 45670 35138 45722
rect 35162 45670 35192 45722
rect 35192 45670 35218 45722
rect 34922 45668 34978 45670
rect 35002 45668 35058 45670
rect 35082 45668 35138 45670
rect 35162 45668 35218 45670
rect 34922 44634 34978 44636
rect 35002 44634 35058 44636
rect 35082 44634 35138 44636
rect 35162 44634 35218 44636
rect 34922 44582 34948 44634
rect 34948 44582 34978 44634
rect 35002 44582 35012 44634
rect 35012 44582 35058 44634
rect 35082 44582 35128 44634
rect 35128 44582 35138 44634
rect 35162 44582 35192 44634
rect 35192 44582 35218 44634
rect 34922 44580 34978 44582
rect 35002 44580 35058 44582
rect 35082 44580 35138 44582
rect 35162 44580 35218 44582
rect 34922 43546 34978 43548
rect 35002 43546 35058 43548
rect 35082 43546 35138 43548
rect 35162 43546 35218 43548
rect 34922 43494 34948 43546
rect 34948 43494 34978 43546
rect 35002 43494 35012 43546
rect 35012 43494 35058 43546
rect 35082 43494 35128 43546
rect 35128 43494 35138 43546
rect 35162 43494 35192 43546
rect 35192 43494 35218 43546
rect 34922 43492 34978 43494
rect 35002 43492 35058 43494
rect 35082 43492 35138 43494
rect 35162 43492 35218 43494
rect 34922 42458 34978 42460
rect 35002 42458 35058 42460
rect 35082 42458 35138 42460
rect 35162 42458 35218 42460
rect 34922 42406 34948 42458
rect 34948 42406 34978 42458
rect 35002 42406 35012 42458
rect 35012 42406 35058 42458
rect 35082 42406 35128 42458
rect 35128 42406 35138 42458
rect 35162 42406 35192 42458
rect 35192 42406 35218 42458
rect 34922 42404 34978 42406
rect 35002 42404 35058 42406
rect 35082 42404 35138 42406
rect 35162 42404 35218 42406
rect 34922 41370 34978 41372
rect 35002 41370 35058 41372
rect 35082 41370 35138 41372
rect 35162 41370 35218 41372
rect 34922 41318 34948 41370
rect 34948 41318 34978 41370
rect 35002 41318 35012 41370
rect 35012 41318 35058 41370
rect 35082 41318 35128 41370
rect 35128 41318 35138 41370
rect 35162 41318 35192 41370
rect 35192 41318 35218 41370
rect 34922 41316 34978 41318
rect 35002 41316 35058 41318
rect 35082 41316 35138 41318
rect 35162 41316 35218 41318
rect 34922 40282 34978 40284
rect 35002 40282 35058 40284
rect 35082 40282 35138 40284
rect 35162 40282 35218 40284
rect 34922 40230 34948 40282
rect 34948 40230 34978 40282
rect 35002 40230 35012 40282
rect 35012 40230 35058 40282
rect 35082 40230 35128 40282
rect 35128 40230 35138 40282
rect 35162 40230 35192 40282
rect 35192 40230 35218 40282
rect 34922 40228 34978 40230
rect 35002 40228 35058 40230
rect 35082 40228 35138 40230
rect 35162 40228 35218 40230
rect 34922 39194 34978 39196
rect 35002 39194 35058 39196
rect 35082 39194 35138 39196
rect 35162 39194 35218 39196
rect 34922 39142 34948 39194
rect 34948 39142 34978 39194
rect 35002 39142 35012 39194
rect 35012 39142 35058 39194
rect 35082 39142 35128 39194
rect 35128 39142 35138 39194
rect 35162 39142 35192 39194
rect 35192 39142 35218 39194
rect 34922 39140 34978 39142
rect 35002 39140 35058 39142
rect 35082 39140 35138 39142
rect 35162 39140 35218 39142
rect 34922 38106 34978 38108
rect 35002 38106 35058 38108
rect 35082 38106 35138 38108
rect 35162 38106 35218 38108
rect 34922 38054 34948 38106
rect 34948 38054 34978 38106
rect 35002 38054 35012 38106
rect 35012 38054 35058 38106
rect 35082 38054 35128 38106
rect 35128 38054 35138 38106
rect 35162 38054 35192 38106
rect 35192 38054 35218 38106
rect 34922 38052 34978 38054
rect 35002 38052 35058 38054
rect 35082 38052 35138 38054
rect 35162 38052 35218 38054
rect 34922 37018 34978 37020
rect 35002 37018 35058 37020
rect 35082 37018 35138 37020
rect 35162 37018 35218 37020
rect 34922 36966 34948 37018
rect 34948 36966 34978 37018
rect 35002 36966 35012 37018
rect 35012 36966 35058 37018
rect 35082 36966 35128 37018
rect 35128 36966 35138 37018
rect 35162 36966 35192 37018
rect 35192 36966 35218 37018
rect 34922 36964 34978 36966
rect 35002 36964 35058 36966
rect 35082 36964 35138 36966
rect 35162 36964 35218 36966
rect 34922 35930 34978 35932
rect 35002 35930 35058 35932
rect 35082 35930 35138 35932
rect 35162 35930 35218 35932
rect 34922 35878 34948 35930
rect 34948 35878 34978 35930
rect 35002 35878 35012 35930
rect 35012 35878 35058 35930
rect 35082 35878 35128 35930
rect 35128 35878 35138 35930
rect 35162 35878 35192 35930
rect 35192 35878 35218 35930
rect 34922 35876 34978 35878
rect 35002 35876 35058 35878
rect 35082 35876 35138 35878
rect 35162 35876 35218 35878
rect 34922 34842 34978 34844
rect 35002 34842 35058 34844
rect 35082 34842 35138 34844
rect 35162 34842 35218 34844
rect 34922 34790 34948 34842
rect 34948 34790 34978 34842
rect 35002 34790 35012 34842
rect 35012 34790 35058 34842
rect 35082 34790 35128 34842
rect 35128 34790 35138 34842
rect 35162 34790 35192 34842
rect 35192 34790 35218 34842
rect 34922 34788 34978 34790
rect 35002 34788 35058 34790
rect 35082 34788 35138 34790
rect 35162 34788 35218 34790
rect 34922 33754 34978 33756
rect 35002 33754 35058 33756
rect 35082 33754 35138 33756
rect 35162 33754 35218 33756
rect 34922 33702 34948 33754
rect 34948 33702 34978 33754
rect 35002 33702 35012 33754
rect 35012 33702 35058 33754
rect 35082 33702 35128 33754
rect 35128 33702 35138 33754
rect 35162 33702 35192 33754
rect 35192 33702 35218 33754
rect 34922 33700 34978 33702
rect 35002 33700 35058 33702
rect 35082 33700 35138 33702
rect 35162 33700 35218 33702
rect 34922 32666 34978 32668
rect 35002 32666 35058 32668
rect 35082 32666 35138 32668
rect 35162 32666 35218 32668
rect 34922 32614 34948 32666
rect 34948 32614 34978 32666
rect 35002 32614 35012 32666
rect 35012 32614 35058 32666
rect 35082 32614 35128 32666
rect 35128 32614 35138 32666
rect 35162 32614 35192 32666
rect 35192 32614 35218 32666
rect 34922 32612 34978 32614
rect 35002 32612 35058 32614
rect 35082 32612 35138 32614
rect 35162 32612 35218 32614
rect 34922 31578 34978 31580
rect 35002 31578 35058 31580
rect 35082 31578 35138 31580
rect 35162 31578 35218 31580
rect 34922 31526 34948 31578
rect 34948 31526 34978 31578
rect 35002 31526 35012 31578
rect 35012 31526 35058 31578
rect 35082 31526 35128 31578
rect 35128 31526 35138 31578
rect 35162 31526 35192 31578
rect 35192 31526 35218 31578
rect 34922 31524 34978 31526
rect 35002 31524 35058 31526
rect 35082 31524 35138 31526
rect 35162 31524 35218 31526
rect 34922 30490 34978 30492
rect 35002 30490 35058 30492
rect 35082 30490 35138 30492
rect 35162 30490 35218 30492
rect 34922 30438 34948 30490
rect 34948 30438 34978 30490
rect 35002 30438 35012 30490
rect 35012 30438 35058 30490
rect 35082 30438 35128 30490
rect 35128 30438 35138 30490
rect 35162 30438 35192 30490
rect 35192 30438 35218 30490
rect 34922 30436 34978 30438
rect 35002 30436 35058 30438
rect 35082 30436 35138 30438
rect 35162 30436 35218 30438
rect 34922 29402 34978 29404
rect 35002 29402 35058 29404
rect 35082 29402 35138 29404
rect 35162 29402 35218 29404
rect 34922 29350 34948 29402
rect 34948 29350 34978 29402
rect 35002 29350 35012 29402
rect 35012 29350 35058 29402
rect 35082 29350 35128 29402
rect 35128 29350 35138 29402
rect 35162 29350 35192 29402
rect 35192 29350 35218 29402
rect 34922 29348 34978 29350
rect 35002 29348 35058 29350
rect 35082 29348 35138 29350
rect 35162 29348 35218 29350
rect 34922 28314 34978 28316
rect 35002 28314 35058 28316
rect 35082 28314 35138 28316
rect 35162 28314 35218 28316
rect 34922 28262 34948 28314
rect 34948 28262 34978 28314
rect 35002 28262 35012 28314
rect 35012 28262 35058 28314
rect 35082 28262 35128 28314
rect 35128 28262 35138 28314
rect 35162 28262 35192 28314
rect 35192 28262 35218 28314
rect 34922 28260 34978 28262
rect 35002 28260 35058 28262
rect 35082 28260 35138 28262
rect 35162 28260 35218 28262
rect 34922 27226 34978 27228
rect 35002 27226 35058 27228
rect 35082 27226 35138 27228
rect 35162 27226 35218 27228
rect 34922 27174 34948 27226
rect 34948 27174 34978 27226
rect 35002 27174 35012 27226
rect 35012 27174 35058 27226
rect 35082 27174 35128 27226
rect 35128 27174 35138 27226
rect 35162 27174 35192 27226
rect 35192 27174 35218 27226
rect 34922 27172 34978 27174
rect 35002 27172 35058 27174
rect 35082 27172 35138 27174
rect 35162 27172 35218 27174
rect 34922 26138 34978 26140
rect 35002 26138 35058 26140
rect 35082 26138 35138 26140
rect 35162 26138 35218 26140
rect 34922 26086 34948 26138
rect 34948 26086 34978 26138
rect 35002 26086 35012 26138
rect 35012 26086 35058 26138
rect 35082 26086 35128 26138
rect 35128 26086 35138 26138
rect 35162 26086 35192 26138
rect 35192 26086 35218 26138
rect 34922 26084 34978 26086
rect 35002 26084 35058 26086
rect 35082 26084 35138 26086
rect 35162 26084 35218 26086
rect 34922 25050 34978 25052
rect 35002 25050 35058 25052
rect 35082 25050 35138 25052
rect 35162 25050 35218 25052
rect 34922 24998 34948 25050
rect 34948 24998 34978 25050
rect 35002 24998 35012 25050
rect 35012 24998 35058 25050
rect 35082 24998 35128 25050
rect 35128 24998 35138 25050
rect 35162 24998 35192 25050
rect 35192 24998 35218 25050
rect 34922 24996 34978 24998
rect 35002 24996 35058 24998
rect 35082 24996 35138 24998
rect 35162 24996 35218 24998
rect 34922 23962 34978 23964
rect 35002 23962 35058 23964
rect 35082 23962 35138 23964
rect 35162 23962 35218 23964
rect 34922 23910 34948 23962
rect 34948 23910 34978 23962
rect 35002 23910 35012 23962
rect 35012 23910 35058 23962
rect 35082 23910 35128 23962
rect 35128 23910 35138 23962
rect 35162 23910 35192 23962
rect 35192 23910 35218 23962
rect 34922 23908 34978 23910
rect 35002 23908 35058 23910
rect 35082 23908 35138 23910
rect 35162 23908 35218 23910
rect 34922 22874 34978 22876
rect 35002 22874 35058 22876
rect 35082 22874 35138 22876
rect 35162 22874 35218 22876
rect 34922 22822 34948 22874
rect 34948 22822 34978 22874
rect 35002 22822 35012 22874
rect 35012 22822 35058 22874
rect 35082 22822 35128 22874
rect 35128 22822 35138 22874
rect 35162 22822 35192 22874
rect 35192 22822 35218 22874
rect 34922 22820 34978 22822
rect 35002 22820 35058 22822
rect 35082 22820 35138 22822
rect 35162 22820 35218 22822
rect 34922 21786 34978 21788
rect 35002 21786 35058 21788
rect 35082 21786 35138 21788
rect 35162 21786 35218 21788
rect 34922 21734 34948 21786
rect 34948 21734 34978 21786
rect 35002 21734 35012 21786
rect 35012 21734 35058 21786
rect 35082 21734 35128 21786
rect 35128 21734 35138 21786
rect 35162 21734 35192 21786
rect 35192 21734 35218 21786
rect 34922 21732 34978 21734
rect 35002 21732 35058 21734
rect 35082 21732 35138 21734
rect 35162 21732 35218 21734
rect 34922 20698 34978 20700
rect 35002 20698 35058 20700
rect 35082 20698 35138 20700
rect 35162 20698 35218 20700
rect 34922 20646 34948 20698
rect 34948 20646 34978 20698
rect 35002 20646 35012 20698
rect 35012 20646 35058 20698
rect 35082 20646 35128 20698
rect 35128 20646 35138 20698
rect 35162 20646 35192 20698
rect 35192 20646 35218 20698
rect 34922 20644 34978 20646
rect 35002 20644 35058 20646
rect 35082 20644 35138 20646
rect 35162 20644 35218 20646
rect 34922 19610 34978 19612
rect 35002 19610 35058 19612
rect 35082 19610 35138 19612
rect 35162 19610 35218 19612
rect 34922 19558 34948 19610
rect 34948 19558 34978 19610
rect 35002 19558 35012 19610
rect 35012 19558 35058 19610
rect 35082 19558 35128 19610
rect 35128 19558 35138 19610
rect 35162 19558 35192 19610
rect 35192 19558 35218 19610
rect 34922 19556 34978 19558
rect 35002 19556 35058 19558
rect 35082 19556 35138 19558
rect 35162 19556 35218 19558
rect 34922 18522 34978 18524
rect 35002 18522 35058 18524
rect 35082 18522 35138 18524
rect 35162 18522 35218 18524
rect 34922 18470 34948 18522
rect 34948 18470 34978 18522
rect 35002 18470 35012 18522
rect 35012 18470 35058 18522
rect 35082 18470 35128 18522
rect 35128 18470 35138 18522
rect 35162 18470 35192 18522
rect 35192 18470 35218 18522
rect 34922 18468 34978 18470
rect 35002 18468 35058 18470
rect 35082 18468 35138 18470
rect 35162 18468 35218 18470
rect 34922 17434 34978 17436
rect 35002 17434 35058 17436
rect 35082 17434 35138 17436
rect 35162 17434 35218 17436
rect 34922 17382 34948 17434
rect 34948 17382 34978 17434
rect 35002 17382 35012 17434
rect 35012 17382 35058 17434
rect 35082 17382 35128 17434
rect 35128 17382 35138 17434
rect 35162 17382 35192 17434
rect 35192 17382 35218 17434
rect 34922 17380 34978 17382
rect 35002 17380 35058 17382
rect 35082 17380 35138 17382
rect 35162 17380 35218 17382
rect 34922 16346 34978 16348
rect 35002 16346 35058 16348
rect 35082 16346 35138 16348
rect 35162 16346 35218 16348
rect 34922 16294 34948 16346
rect 34948 16294 34978 16346
rect 35002 16294 35012 16346
rect 35012 16294 35058 16346
rect 35082 16294 35128 16346
rect 35128 16294 35138 16346
rect 35162 16294 35192 16346
rect 35192 16294 35218 16346
rect 34922 16292 34978 16294
rect 35002 16292 35058 16294
rect 35082 16292 35138 16294
rect 35162 16292 35218 16294
rect 34040 3712 34096 3768
rect 34500 3168 34556 3224
rect 34500 2896 34556 2952
rect 34922 15258 34978 15260
rect 35002 15258 35058 15260
rect 35082 15258 35138 15260
rect 35162 15258 35218 15260
rect 34922 15206 34948 15258
rect 34948 15206 34978 15258
rect 35002 15206 35012 15258
rect 35012 15206 35058 15258
rect 35082 15206 35128 15258
rect 35128 15206 35138 15258
rect 35162 15206 35192 15258
rect 35192 15206 35218 15258
rect 34922 15204 34978 15206
rect 35002 15204 35058 15206
rect 35082 15204 35138 15206
rect 35162 15204 35218 15206
rect 34922 14170 34978 14172
rect 35002 14170 35058 14172
rect 35082 14170 35138 14172
rect 35162 14170 35218 14172
rect 34922 14118 34948 14170
rect 34948 14118 34978 14170
rect 35002 14118 35012 14170
rect 35012 14118 35058 14170
rect 35082 14118 35128 14170
rect 35128 14118 35138 14170
rect 35162 14118 35192 14170
rect 35192 14118 35218 14170
rect 34922 14116 34978 14118
rect 35002 14116 35058 14118
rect 35082 14116 35138 14118
rect 35162 14116 35218 14118
rect 34922 13082 34978 13084
rect 35002 13082 35058 13084
rect 35082 13082 35138 13084
rect 35162 13082 35218 13084
rect 34922 13030 34948 13082
rect 34948 13030 34978 13082
rect 35002 13030 35012 13082
rect 35012 13030 35058 13082
rect 35082 13030 35128 13082
rect 35128 13030 35138 13082
rect 35162 13030 35192 13082
rect 35192 13030 35218 13082
rect 34922 13028 34978 13030
rect 35002 13028 35058 13030
rect 35082 13028 35138 13030
rect 35162 13028 35218 13030
rect 34922 11994 34978 11996
rect 35002 11994 35058 11996
rect 35082 11994 35138 11996
rect 35162 11994 35218 11996
rect 34922 11942 34948 11994
rect 34948 11942 34978 11994
rect 35002 11942 35012 11994
rect 35012 11942 35058 11994
rect 35082 11942 35128 11994
rect 35128 11942 35138 11994
rect 35162 11942 35192 11994
rect 35192 11942 35218 11994
rect 34922 11940 34978 11942
rect 35002 11940 35058 11942
rect 35082 11940 35138 11942
rect 35162 11940 35218 11942
rect 34922 10906 34978 10908
rect 35002 10906 35058 10908
rect 35082 10906 35138 10908
rect 35162 10906 35218 10908
rect 34922 10854 34948 10906
rect 34948 10854 34978 10906
rect 35002 10854 35012 10906
rect 35012 10854 35058 10906
rect 35082 10854 35128 10906
rect 35128 10854 35138 10906
rect 35162 10854 35192 10906
rect 35192 10854 35218 10906
rect 34922 10852 34978 10854
rect 35002 10852 35058 10854
rect 35082 10852 35138 10854
rect 35162 10852 35218 10854
rect 34922 9818 34978 9820
rect 35002 9818 35058 9820
rect 35082 9818 35138 9820
rect 35162 9818 35218 9820
rect 34922 9766 34948 9818
rect 34948 9766 34978 9818
rect 35002 9766 35012 9818
rect 35012 9766 35058 9818
rect 35082 9766 35128 9818
rect 35128 9766 35138 9818
rect 35162 9766 35192 9818
rect 35192 9766 35218 9818
rect 34922 9764 34978 9766
rect 35002 9764 35058 9766
rect 35082 9764 35138 9766
rect 35162 9764 35218 9766
rect 34922 8730 34978 8732
rect 35002 8730 35058 8732
rect 35082 8730 35138 8732
rect 35162 8730 35218 8732
rect 34922 8678 34948 8730
rect 34948 8678 34978 8730
rect 35002 8678 35012 8730
rect 35012 8678 35058 8730
rect 35082 8678 35128 8730
rect 35128 8678 35138 8730
rect 35162 8678 35192 8730
rect 35192 8678 35218 8730
rect 34922 8676 34978 8678
rect 35002 8676 35058 8678
rect 35082 8676 35138 8678
rect 35162 8676 35218 8678
rect 34922 7642 34978 7644
rect 35002 7642 35058 7644
rect 35082 7642 35138 7644
rect 35162 7642 35218 7644
rect 34922 7590 34948 7642
rect 34948 7590 34978 7642
rect 35002 7590 35012 7642
rect 35012 7590 35058 7642
rect 35082 7590 35128 7642
rect 35128 7590 35138 7642
rect 35162 7590 35192 7642
rect 35192 7590 35218 7642
rect 34922 7588 34978 7590
rect 35002 7588 35058 7590
rect 35082 7588 35138 7590
rect 35162 7588 35218 7590
rect 34922 6554 34978 6556
rect 35002 6554 35058 6556
rect 35082 6554 35138 6556
rect 35162 6554 35218 6556
rect 34922 6502 34948 6554
rect 34948 6502 34978 6554
rect 35002 6502 35012 6554
rect 35012 6502 35058 6554
rect 35082 6502 35128 6554
rect 35128 6502 35138 6554
rect 35162 6502 35192 6554
rect 35192 6502 35218 6554
rect 34922 6500 34978 6502
rect 35002 6500 35058 6502
rect 35082 6500 35138 6502
rect 35162 6500 35218 6502
rect 34922 5466 34978 5468
rect 35002 5466 35058 5468
rect 35082 5466 35138 5468
rect 35162 5466 35218 5468
rect 34922 5414 34948 5466
rect 34948 5414 34978 5466
rect 35002 5414 35012 5466
rect 35012 5414 35058 5466
rect 35082 5414 35128 5466
rect 35128 5414 35138 5466
rect 35162 5414 35192 5466
rect 35192 5414 35218 5466
rect 34922 5412 34978 5414
rect 35002 5412 35058 5414
rect 35082 5412 35138 5414
rect 35162 5412 35218 5414
rect 34922 4378 34978 4380
rect 35002 4378 35058 4380
rect 35082 4378 35138 4380
rect 35162 4378 35218 4380
rect 34922 4326 34948 4378
rect 34948 4326 34978 4378
rect 35002 4326 35012 4378
rect 35012 4326 35058 4378
rect 35082 4326 35128 4378
rect 35128 4326 35138 4378
rect 35162 4326 35192 4378
rect 35192 4326 35218 4378
rect 34922 4324 34978 4326
rect 35002 4324 35058 4326
rect 35082 4324 35138 4326
rect 35162 4324 35218 4326
rect 34922 3290 34978 3292
rect 35002 3290 35058 3292
rect 35082 3290 35138 3292
rect 35162 3290 35218 3292
rect 34922 3238 34948 3290
rect 34948 3238 34978 3290
rect 35002 3238 35012 3290
rect 35012 3238 35058 3290
rect 35082 3238 35128 3290
rect 35128 3238 35138 3290
rect 35162 3238 35192 3290
rect 35192 3238 35218 3290
rect 34922 3236 34978 3238
rect 35002 3236 35058 3238
rect 35082 3236 35138 3238
rect 35162 3236 35218 3238
rect 35420 2896 35476 2952
rect 34922 2202 34978 2204
rect 35002 2202 35058 2204
rect 35082 2202 35138 2204
rect 35162 2202 35218 2204
rect 34922 2150 34948 2202
rect 34948 2150 34978 2202
rect 35002 2150 35012 2202
rect 35012 2150 35058 2202
rect 35082 2150 35128 2202
rect 35128 2150 35138 2202
rect 35162 2150 35192 2202
rect 35192 2150 35218 2202
rect 34922 2148 34978 2150
rect 35002 2148 35058 2150
rect 35082 2148 35138 2150
rect 35162 2148 35218 2150
rect 37352 16496 37408 16552
rect 37628 2760 37684 2816
rect 40204 56380 40206 56400
rect 40206 56380 40258 56400
rect 40258 56380 40260 56400
rect 40204 56344 40260 56380
rect 41124 56364 41180 56400
rect 41124 56344 41126 56364
rect 41126 56344 41178 56364
rect 41178 56344 41180 56364
rect 41308 56208 41364 56264
rect 41492 56344 41548 56400
rect 38824 44104 38880 44160
rect 38732 16632 38788 16688
rect 38640 2896 38696 2952
rect 39008 26288 39064 26344
rect 41308 55412 41364 55448
rect 41308 55392 41310 55412
rect 41310 55392 41362 55412
rect 41362 55392 41364 55412
rect 42044 3032 42100 3088
rect 41124 2896 41180 2952
rect 43516 3984 43572 4040
rect 45448 55392 45504 55448
rect 50282 57146 50338 57148
rect 50362 57146 50418 57148
rect 50442 57146 50498 57148
rect 50522 57146 50578 57148
rect 50282 57094 50308 57146
rect 50308 57094 50338 57146
rect 50362 57094 50372 57146
rect 50372 57094 50418 57146
rect 50442 57094 50488 57146
rect 50488 57094 50498 57146
rect 50522 57094 50552 57146
rect 50552 57094 50578 57146
rect 50282 57092 50338 57094
rect 50362 57092 50418 57094
rect 50442 57092 50498 57094
rect 50522 57092 50578 57094
rect 51244 57976 51300 58032
rect 50282 56058 50338 56060
rect 50362 56058 50418 56060
rect 50442 56058 50498 56060
rect 50522 56058 50578 56060
rect 50282 56006 50308 56058
rect 50308 56006 50338 56058
rect 50362 56006 50372 56058
rect 50372 56006 50418 56058
rect 50442 56006 50488 56058
rect 50488 56006 50498 56058
rect 50522 56006 50552 56058
rect 50552 56006 50578 56058
rect 50282 56004 50338 56006
rect 50362 56004 50418 56006
rect 50442 56004 50498 56006
rect 50522 56004 50578 56006
rect 45540 53760 45596 53816
rect 45724 53760 45780 53816
rect 44620 3712 44676 3768
rect 45540 34448 45596 34504
rect 45724 34448 45780 34504
rect 45356 24792 45412 24848
rect 45724 24828 45726 24848
rect 45726 24828 45778 24848
rect 45778 24828 45780 24848
rect 45724 24792 45780 24828
rect 47196 3576 47252 3632
rect 48300 19216 48356 19272
rect 48392 19080 48448 19136
rect 49220 9560 49276 9616
rect 48392 3304 48448 3360
rect 50282 54970 50338 54972
rect 50362 54970 50418 54972
rect 50442 54970 50498 54972
rect 50522 54970 50578 54972
rect 50282 54918 50308 54970
rect 50308 54918 50338 54970
rect 50362 54918 50372 54970
rect 50372 54918 50418 54970
rect 50442 54918 50488 54970
rect 50488 54918 50498 54970
rect 50522 54918 50552 54970
rect 50552 54918 50578 54970
rect 50282 54916 50338 54918
rect 50362 54916 50418 54918
rect 50442 54916 50498 54918
rect 50522 54916 50578 54918
rect 50282 53882 50338 53884
rect 50362 53882 50418 53884
rect 50442 53882 50498 53884
rect 50522 53882 50578 53884
rect 50282 53830 50308 53882
rect 50308 53830 50338 53882
rect 50362 53830 50372 53882
rect 50372 53830 50418 53882
rect 50442 53830 50488 53882
rect 50488 53830 50498 53882
rect 50522 53830 50552 53882
rect 50552 53830 50578 53882
rect 50282 53828 50338 53830
rect 50362 53828 50418 53830
rect 50442 53828 50498 53830
rect 50522 53828 50578 53830
rect 52256 57976 52312 58032
rect 50282 52794 50338 52796
rect 50362 52794 50418 52796
rect 50442 52794 50498 52796
rect 50522 52794 50578 52796
rect 50282 52742 50308 52794
rect 50308 52742 50338 52794
rect 50362 52742 50372 52794
rect 50372 52742 50418 52794
rect 50442 52742 50488 52794
rect 50488 52742 50498 52794
rect 50522 52742 50552 52794
rect 50552 52742 50578 52794
rect 50282 52740 50338 52742
rect 50362 52740 50418 52742
rect 50442 52740 50498 52742
rect 50522 52740 50578 52742
rect 50282 51706 50338 51708
rect 50362 51706 50418 51708
rect 50442 51706 50498 51708
rect 50522 51706 50578 51708
rect 50282 51654 50308 51706
rect 50308 51654 50338 51706
rect 50362 51654 50372 51706
rect 50372 51654 50418 51706
rect 50442 51654 50488 51706
rect 50488 51654 50498 51706
rect 50522 51654 50552 51706
rect 50552 51654 50578 51706
rect 50282 51652 50338 51654
rect 50362 51652 50418 51654
rect 50442 51652 50498 51654
rect 50522 51652 50578 51654
rect 50282 50618 50338 50620
rect 50362 50618 50418 50620
rect 50442 50618 50498 50620
rect 50522 50618 50578 50620
rect 50282 50566 50308 50618
rect 50308 50566 50338 50618
rect 50362 50566 50372 50618
rect 50372 50566 50418 50618
rect 50442 50566 50488 50618
rect 50488 50566 50498 50618
rect 50522 50566 50552 50618
rect 50552 50566 50578 50618
rect 50282 50564 50338 50566
rect 50362 50564 50418 50566
rect 50442 50564 50498 50566
rect 50522 50564 50578 50566
rect 50282 49530 50338 49532
rect 50362 49530 50418 49532
rect 50442 49530 50498 49532
rect 50522 49530 50578 49532
rect 50282 49478 50308 49530
rect 50308 49478 50338 49530
rect 50362 49478 50372 49530
rect 50372 49478 50418 49530
rect 50442 49478 50488 49530
rect 50488 49478 50498 49530
rect 50522 49478 50552 49530
rect 50552 49478 50578 49530
rect 50282 49476 50338 49478
rect 50362 49476 50418 49478
rect 50442 49476 50498 49478
rect 50522 49476 50578 49478
rect 50282 48442 50338 48444
rect 50362 48442 50418 48444
rect 50442 48442 50498 48444
rect 50522 48442 50578 48444
rect 50282 48390 50308 48442
rect 50308 48390 50338 48442
rect 50362 48390 50372 48442
rect 50372 48390 50418 48442
rect 50442 48390 50488 48442
rect 50488 48390 50498 48442
rect 50522 48390 50552 48442
rect 50552 48390 50578 48442
rect 50282 48388 50338 48390
rect 50362 48388 50418 48390
rect 50442 48388 50498 48390
rect 50522 48388 50578 48390
rect 50282 47354 50338 47356
rect 50362 47354 50418 47356
rect 50442 47354 50498 47356
rect 50522 47354 50578 47356
rect 50282 47302 50308 47354
rect 50308 47302 50338 47354
rect 50362 47302 50372 47354
rect 50372 47302 50418 47354
rect 50442 47302 50488 47354
rect 50488 47302 50498 47354
rect 50522 47302 50552 47354
rect 50552 47302 50578 47354
rect 50282 47300 50338 47302
rect 50362 47300 50418 47302
rect 50442 47300 50498 47302
rect 50522 47300 50578 47302
rect 50282 46266 50338 46268
rect 50362 46266 50418 46268
rect 50442 46266 50498 46268
rect 50522 46266 50578 46268
rect 50282 46214 50308 46266
rect 50308 46214 50338 46266
rect 50362 46214 50372 46266
rect 50372 46214 50418 46266
rect 50442 46214 50488 46266
rect 50488 46214 50498 46266
rect 50522 46214 50552 46266
rect 50552 46214 50578 46266
rect 50282 46212 50338 46214
rect 50362 46212 50418 46214
rect 50442 46212 50498 46214
rect 50522 46212 50578 46214
rect 50282 45178 50338 45180
rect 50362 45178 50418 45180
rect 50442 45178 50498 45180
rect 50522 45178 50578 45180
rect 50282 45126 50308 45178
rect 50308 45126 50338 45178
rect 50362 45126 50372 45178
rect 50372 45126 50418 45178
rect 50442 45126 50488 45178
rect 50488 45126 50498 45178
rect 50522 45126 50552 45178
rect 50552 45126 50578 45178
rect 50282 45124 50338 45126
rect 50362 45124 50418 45126
rect 50442 45124 50498 45126
rect 50522 45124 50578 45126
rect 50282 44090 50338 44092
rect 50362 44090 50418 44092
rect 50442 44090 50498 44092
rect 50522 44090 50578 44092
rect 50282 44038 50308 44090
rect 50308 44038 50338 44090
rect 50362 44038 50372 44090
rect 50372 44038 50418 44090
rect 50442 44038 50488 44090
rect 50488 44038 50498 44090
rect 50522 44038 50552 44090
rect 50552 44038 50578 44090
rect 50282 44036 50338 44038
rect 50362 44036 50418 44038
rect 50442 44036 50498 44038
rect 50522 44036 50578 44038
rect 50282 43002 50338 43004
rect 50362 43002 50418 43004
rect 50442 43002 50498 43004
rect 50522 43002 50578 43004
rect 50282 42950 50308 43002
rect 50308 42950 50338 43002
rect 50362 42950 50372 43002
rect 50372 42950 50418 43002
rect 50442 42950 50488 43002
rect 50488 42950 50498 43002
rect 50522 42950 50552 43002
rect 50552 42950 50578 43002
rect 50282 42948 50338 42950
rect 50362 42948 50418 42950
rect 50442 42948 50498 42950
rect 50522 42948 50578 42950
rect 50282 41914 50338 41916
rect 50362 41914 50418 41916
rect 50442 41914 50498 41916
rect 50522 41914 50578 41916
rect 50282 41862 50308 41914
rect 50308 41862 50338 41914
rect 50362 41862 50372 41914
rect 50372 41862 50418 41914
rect 50442 41862 50488 41914
rect 50488 41862 50498 41914
rect 50522 41862 50552 41914
rect 50552 41862 50578 41914
rect 50282 41860 50338 41862
rect 50362 41860 50418 41862
rect 50442 41860 50498 41862
rect 50522 41860 50578 41862
rect 50282 40826 50338 40828
rect 50362 40826 50418 40828
rect 50442 40826 50498 40828
rect 50522 40826 50578 40828
rect 50282 40774 50308 40826
rect 50308 40774 50338 40826
rect 50362 40774 50372 40826
rect 50372 40774 50418 40826
rect 50442 40774 50488 40826
rect 50488 40774 50498 40826
rect 50522 40774 50552 40826
rect 50552 40774 50578 40826
rect 50282 40772 50338 40774
rect 50362 40772 50418 40774
rect 50442 40772 50498 40774
rect 50522 40772 50578 40774
rect 50282 39738 50338 39740
rect 50362 39738 50418 39740
rect 50442 39738 50498 39740
rect 50522 39738 50578 39740
rect 50282 39686 50308 39738
rect 50308 39686 50338 39738
rect 50362 39686 50372 39738
rect 50372 39686 50418 39738
rect 50442 39686 50488 39738
rect 50488 39686 50498 39738
rect 50522 39686 50552 39738
rect 50552 39686 50578 39738
rect 50282 39684 50338 39686
rect 50362 39684 50418 39686
rect 50442 39684 50498 39686
rect 50522 39684 50578 39686
rect 50282 38650 50338 38652
rect 50362 38650 50418 38652
rect 50442 38650 50498 38652
rect 50522 38650 50578 38652
rect 50282 38598 50308 38650
rect 50308 38598 50338 38650
rect 50362 38598 50372 38650
rect 50372 38598 50418 38650
rect 50442 38598 50488 38650
rect 50488 38598 50498 38650
rect 50522 38598 50552 38650
rect 50552 38598 50578 38650
rect 50282 38596 50338 38598
rect 50362 38596 50418 38598
rect 50442 38596 50498 38598
rect 50522 38596 50578 38598
rect 50282 37562 50338 37564
rect 50362 37562 50418 37564
rect 50442 37562 50498 37564
rect 50522 37562 50578 37564
rect 50282 37510 50308 37562
rect 50308 37510 50338 37562
rect 50362 37510 50372 37562
rect 50372 37510 50418 37562
rect 50442 37510 50488 37562
rect 50488 37510 50498 37562
rect 50522 37510 50552 37562
rect 50552 37510 50578 37562
rect 50282 37508 50338 37510
rect 50362 37508 50418 37510
rect 50442 37508 50498 37510
rect 50522 37508 50578 37510
rect 50282 36474 50338 36476
rect 50362 36474 50418 36476
rect 50442 36474 50498 36476
rect 50522 36474 50578 36476
rect 50282 36422 50308 36474
rect 50308 36422 50338 36474
rect 50362 36422 50372 36474
rect 50372 36422 50418 36474
rect 50442 36422 50488 36474
rect 50488 36422 50498 36474
rect 50522 36422 50552 36474
rect 50552 36422 50578 36474
rect 50282 36420 50338 36422
rect 50362 36420 50418 36422
rect 50442 36420 50498 36422
rect 50522 36420 50578 36422
rect 50282 35386 50338 35388
rect 50362 35386 50418 35388
rect 50442 35386 50498 35388
rect 50522 35386 50578 35388
rect 50282 35334 50308 35386
rect 50308 35334 50338 35386
rect 50362 35334 50372 35386
rect 50372 35334 50418 35386
rect 50442 35334 50488 35386
rect 50488 35334 50498 35386
rect 50522 35334 50552 35386
rect 50552 35334 50578 35386
rect 50282 35332 50338 35334
rect 50362 35332 50418 35334
rect 50442 35332 50498 35334
rect 50522 35332 50578 35334
rect 50282 34298 50338 34300
rect 50362 34298 50418 34300
rect 50442 34298 50498 34300
rect 50522 34298 50578 34300
rect 50282 34246 50308 34298
rect 50308 34246 50338 34298
rect 50362 34246 50372 34298
rect 50372 34246 50418 34298
rect 50442 34246 50488 34298
rect 50488 34246 50498 34298
rect 50522 34246 50552 34298
rect 50552 34246 50578 34298
rect 50282 34244 50338 34246
rect 50362 34244 50418 34246
rect 50442 34244 50498 34246
rect 50522 34244 50578 34246
rect 50282 33210 50338 33212
rect 50362 33210 50418 33212
rect 50442 33210 50498 33212
rect 50522 33210 50578 33212
rect 50282 33158 50308 33210
rect 50308 33158 50338 33210
rect 50362 33158 50372 33210
rect 50372 33158 50418 33210
rect 50442 33158 50488 33210
rect 50488 33158 50498 33210
rect 50522 33158 50552 33210
rect 50552 33158 50578 33210
rect 50282 33156 50338 33158
rect 50362 33156 50418 33158
rect 50442 33156 50498 33158
rect 50522 33156 50578 33158
rect 50282 32122 50338 32124
rect 50362 32122 50418 32124
rect 50442 32122 50498 32124
rect 50522 32122 50578 32124
rect 50282 32070 50308 32122
rect 50308 32070 50338 32122
rect 50362 32070 50372 32122
rect 50372 32070 50418 32122
rect 50442 32070 50488 32122
rect 50488 32070 50498 32122
rect 50522 32070 50552 32122
rect 50552 32070 50578 32122
rect 50282 32068 50338 32070
rect 50362 32068 50418 32070
rect 50442 32068 50498 32070
rect 50522 32068 50578 32070
rect 50282 31034 50338 31036
rect 50362 31034 50418 31036
rect 50442 31034 50498 31036
rect 50522 31034 50578 31036
rect 50282 30982 50308 31034
rect 50308 30982 50338 31034
rect 50362 30982 50372 31034
rect 50372 30982 50418 31034
rect 50442 30982 50488 31034
rect 50488 30982 50498 31034
rect 50522 30982 50552 31034
rect 50552 30982 50578 31034
rect 50282 30980 50338 30982
rect 50362 30980 50418 30982
rect 50442 30980 50498 30982
rect 50522 30980 50578 30982
rect 50282 29946 50338 29948
rect 50362 29946 50418 29948
rect 50442 29946 50498 29948
rect 50522 29946 50578 29948
rect 50282 29894 50308 29946
rect 50308 29894 50338 29946
rect 50362 29894 50372 29946
rect 50372 29894 50418 29946
rect 50442 29894 50488 29946
rect 50488 29894 50498 29946
rect 50522 29894 50552 29946
rect 50552 29894 50578 29946
rect 50282 29892 50338 29894
rect 50362 29892 50418 29894
rect 50442 29892 50498 29894
rect 50522 29892 50578 29894
rect 50282 28858 50338 28860
rect 50362 28858 50418 28860
rect 50442 28858 50498 28860
rect 50522 28858 50578 28860
rect 50282 28806 50308 28858
rect 50308 28806 50338 28858
rect 50362 28806 50372 28858
rect 50372 28806 50418 28858
rect 50442 28806 50488 28858
rect 50488 28806 50498 28858
rect 50522 28806 50552 28858
rect 50552 28806 50578 28858
rect 50282 28804 50338 28806
rect 50362 28804 50418 28806
rect 50442 28804 50498 28806
rect 50522 28804 50578 28806
rect 50282 27770 50338 27772
rect 50362 27770 50418 27772
rect 50442 27770 50498 27772
rect 50522 27770 50578 27772
rect 50282 27718 50308 27770
rect 50308 27718 50338 27770
rect 50362 27718 50372 27770
rect 50372 27718 50418 27770
rect 50442 27718 50488 27770
rect 50488 27718 50498 27770
rect 50522 27718 50552 27770
rect 50552 27718 50578 27770
rect 50282 27716 50338 27718
rect 50362 27716 50418 27718
rect 50442 27716 50498 27718
rect 50522 27716 50578 27718
rect 50282 26682 50338 26684
rect 50362 26682 50418 26684
rect 50442 26682 50498 26684
rect 50522 26682 50578 26684
rect 50282 26630 50308 26682
rect 50308 26630 50338 26682
rect 50362 26630 50372 26682
rect 50372 26630 50418 26682
rect 50442 26630 50488 26682
rect 50488 26630 50498 26682
rect 50522 26630 50552 26682
rect 50552 26630 50578 26682
rect 50282 26628 50338 26630
rect 50362 26628 50418 26630
rect 50442 26628 50498 26630
rect 50522 26628 50578 26630
rect 50282 25594 50338 25596
rect 50362 25594 50418 25596
rect 50442 25594 50498 25596
rect 50522 25594 50578 25596
rect 50282 25542 50308 25594
rect 50308 25542 50338 25594
rect 50362 25542 50372 25594
rect 50372 25542 50418 25594
rect 50442 25542 50488 25594
rect 50488 25542 50498 25594
rect 50522 25542 50552 25594
rect 50552 25542 50578 25594
rect 50282 25540 50338 25542
rect 50362 25540 50418 25542
rect 50442 25540 50498 25542
rect 50522 25540 50578 25542
rect 50282 24506 50338 24508
rect 50362 24506 50418 24508
rect 50442 24506 50498 24508
rect 50522 24506 50578 24508
rect 50282 24454 50308 24506
rect 50308 24454 50338 24506
rect 50362 24454 50372 24506
rect 50372 24454 50418 24506
rect 50442 24454 50488 24506
rect 50488 24454 50498 24506
rect 50522 24454 50552 24506
rect 50552 24454 50578 24506
rect 50282 24452 50338 24454
rect 50362 24452 50418 24454
rect 50442 24452 50498 24454
rect 50522 24452 50578 24454
rect 50282 23418 50338 23420
rect 50362 23418 50418 23420
rect 50442 23418 50498 23420
rect 50522 23418 50578 23420
rect 50282 23366 50308 23418
rect 50308 23366 50338 23418
rect 50362 23366 50372 23418
rect 50372 23366 50418 23418
rect 50442 23366 50488 23418
rect 50488 23366 50498 23418
rect 50522 23366 50552 23418
rect 50552 23366 50578 23418
rect 50282 23364 50338 23366
rect 50362 23364 50418 23366
rect 50442 23364 50498 23366
rect 50522 23364 50578 23366
rect 50282 22330 50338 22332
rect 50362 22330 50418 22332
rect 50442 22330 50498 22332
rect 50522 22330 50578 22332
rect 50282 22278 50308 22330
rect 50308 22278 50338 22330
rect 50362 22278 50372 22330
rect 50372 22278 50418 22330
rect 50442 22278 50488 22330
rect 50488 22278 50498 22330
rect 50522 22278 50552 22330
rect 50552 22278 50578 22330
rect 50282 22276 50338 22278
rect 50362 22276 50418 22278
rect 50442 22276 50498 22278
rect 50522 22276 50578 22278
rect 50282 21242 50338 21244
rect 50362 21242 50418 21244
rect 50442 21242 50498 21244
rect 50522 21242 50578 21244
rect 50282 21190 50308 21242
rect 50308 21190 50338 21242
rect 50362 21190 50372 21242
rect 50372 21190 50418 21242
rect 50442 21190 50488 21242
rect 50488 21190 50498 21242
rect 50522 21190 50552 21242
rect 50552 21190 50578 21242
rect 50282 21188 50338 21190
rect 50362 21188 50418 21190
rect 50442 21188 50498 21190
rect 50522 21188 50578 21190
rect 50282 20154 50338 20156
rect 50362 20154 50418 20156
rect 50442 20154 50498 20156
rect 50522 20154 50578 20156
rect 50282 20102 50308 20154
rect 50308 20102 50338 20154
rect 50362 20102 50372 20154
rect 50372 20102 50418 20154
rect 50442 20102 50488 20154
rect 50488 20102 50498 20154
rect 50522 20102 50552 20154
rect 50552 20102 50578 20154
rect 50282 20100 50338 20102
rect 50362 20100 50418 20102
rect 50442 20100 50498 20102
rect 50522 20100 50578 20102
rect 50282 19066 50338 19068
rect 50362 19066 50418 19068
rect 50442 19066 50498 19068
rect 50522 19066 50578 19068
rect 50282 19014 50308 19066
rect 50308 19014 50338 19066
rect 50362 19014 50372 19066
rect 50372 19014 50418 19066
rect 50442 19014 50488 19066
rect 50488 19014 50498 19066
rect 50522 19014 50552 19066
rect 50552 19014 50578 19066
rect 50282 19012 50338 19014
rect 50362 19012 50418 19014
rect 50442 19012 50498 19014
rect 50522 19012 50578 19014
rect 50282 17978 50338 17980
rect 50362 17978 50418 17980
rect 50442 17978 50498 17980
rect 50522 17978 50578 17980
rect 50282 17926 50308 17978
rect 50308 17926 50338 17978
rect 50362 17926 50372 17978
rect 50372 17926 50418 17978
rect 50442 17926 50488 17978
rect 50488 17926 50498 17978
rect 50522 17926 50552 17978
rect 50552 17926 50578 17978
rect 50282 17924 50338 17926
rect 50362 17924 50418 17926
rect 50442 17924 50498 17926
rect 50522 17924 50578 17926
rect 50282 16890 50338 16892
rect 50362 16890 50418 16892
rect 50442 16890 50498 16892
rect 50522 16890 50578 16892
rect 50282 16838 50308 16890
rect 50308 16838 50338 16890
rect 50362 16838 50372 16890
rect 50372 16838 50418 16890
rect 50442 16838 50488 16890
rect 50488 16838 50498 16890
rect 50522 16838 50552 16890
rect 50552 16838 50578 16890
rect 50282 16836 50338 16838
rect 50362 16836 50418 16838
rect 50442 16836 50498 16838
rect 50522 16836 50578 16838
rect 50282 15802 50338 15804
rect 50362 15802 50418 15804
rect 50442 15802 50498 15804
rect 50522 15802 50578 15804
rect 50282 15750 50308 15802
rect 50308 15750 50338 15802
rect 50362 15750 50372 15802
rect 50372 15750 50418 15802
rect 50442 15750 50488 15802
rect 50488 15750 50498 15802
rect 50522 15750 50552 15802
rect 50552 15750 50578 15802
rect 50282 15748 50338 15750
rect 50362 15748 50418 15750
rect 50442 15748 50498 15750
rect 50522 15748 50578 15750
rect 50282 14714 50338 14716
rect 50362 14714 50418 14716
rect 50442 14714 50498 14716
rect 50522 14714 50578 14716
rect 50282 14662 50308 14714
rect 50308 14662 50338 14714
rect 50362 14662 50372 14714
rect 50372 14662 50418 14714
rect 50442 14662 50488 14714
rect 50488 14662 50498 14714
rect 50522 14662 50552 14714
rect 50552 14662 50578 14714
rect 50282 14660 50338 14662
rect 50362 14660 50418 14662
rect 50442 14660 50498 14662
rect 50522 14660 50578 14662
rect 50282 13626 50338 13628
rect 50362 13626 50418 13628
rect 50442 13626 50498 13628
rect 50522 13626 50578 13628
rect 50282 13574 50308 13626
rect 50308 13574 50338 13626
rect 50362 13574 50372 13626
rect 50372 13574 50418 13626
rect 50442 13574 50488 13626
rect 50488 13574 50498 13626
rect 50522 13574 50552 13626
rect 50552 13574 50578 13626
rect 50282 13572 50338 13574
rect 50362 13572 50418 13574
rect 50442 13572 50498 13574
rect 50522 13572 50578 13574
rect 50282 12538 50338 12540
rect 50362 12538 50418 12540
rect 50442 12538 50498 12540
rect 50522 12538 50578 12540
rect 50282 12486 50308 12538
rect 50308 12486 50338 12538
rect 50362 12486 50372 12538
rect 50372 12486 50418 12538
rect 50442 12486 50488 12538
rect 50488 12486 50498 12538
rect 50522 12486 50552 12538
rect 50552 12486 50578 12538
rect 50282 12484 50338 12486
rect 50362 12484 50418 12486
rect 50442 12484 50498 12486
rect 50522 12484 50578 12486
rect 50282 11450 50338 11452
rect 50362 11450 50418 11452
rect 50442 11450 50498 11452
rect 50522 11450 50578 11452
rect 50282 11398 50308 11450
rect 50308 11398 50338 11450
rect 50362 11398 50372 11450
rect 50372 11398 50418 11450
rect 50442 11398 50488 11450
rect 50488 11398 50498 11450
rect 50522 11398 50552 11450
rect 50552 11398 50578 11450
rect 50282 11396 50338 11398
rect 50362 11396 50418 11398
rect 50442 11396 50498 11398
rect 50522 11396 50578 11398
rect 50282 10362 50338 10364
rect 50362 10362 50418 10364
rect 50442 10362 50498 10364
rect 50522 10362 50578 10364
rect 50282 10310 50308 10362
rect 50308 10310 50338 10362
rect 50362 10310 50372 10362
rect 50372 10310 50418 10362
rect 50442 10310 50488 10362
rect 50488 10310 50498 10362
rect 50522 10310 50552 10362
rect 50552 10310 50578 10362
rect 50282 10308 50338 10310
rect 50362 10308 50418 10310
rect 50442 10308 50498 10310
rect 50522 10308 50578 10310
rect 50282 9274 50338 9276
rect 50362 9274 50418 9276
rect 50442 9274 50498 9276
rect 50522 9274 50578 9276
rect 50282 9222 50308 9274
rect 50308 9222 50338 9274
rect 50362 9222 50372 9274
rect 50372 9222 50418 9274
rect 50442 9222 50488 9274
rect 50488 9222 50498 9274
rect 50522 9222 50552 9274
rect 50552 9222 50578 9274
rect 50282 9220 50338 9222
rect 50362 9220 50418 9222
rect 50442 9220 50498 9222
rect 50522 9220 50578 9222
rect 50282 8186 50338 8188
rect 50362 8186 50418 8188
rect 50442 8186 50498 8188
rect 50522 8186 50578 8188
rect 50282 8134 50308 8186
rect 50308 8134 50338 8186
rect 50362 8134 50372 8186
rect 50372 8134 50418 8186
rect 50442 8134 50488 8186
rect 50488 8134 50498 8186
rect 50522 8134 50552 8186
rect 50552 8134 50578 8186
rect 50282 8132 50338 8134
rect 50362 8132 50418 8134
rect 50442 8132 50498 8134
rect 50522 8132 50578 8134
rect 50282 7098 50338 7100
rect 50362 7098 50418 7100
rect 50442 7098 50498 7100
rect 50522 7098 50578 7100
rect 50282 7046 50308 7098
rect 50308 7046 50338 7098
rect 50362 7046 50372 7098
rect 50372 7046 50418 7098
rect 50442 7046 50488 7098
rect 50488 7046 50498 7098
rect 50522 7046 50552 7098
rect 50552 7046 50578 7098
rect 50282 7044 50338 7046
rect 50362 7044 50418 7046
rect 50442 7044 50498 7046
rect 50522 7044 50578 7046
rect 50282 6010 50338 6012
rect 50362 6010 50418 6012
rect 50442 6010 50498 6012
rect 50522 6010 50578 6012
rect 50282 5958 50308 6010
rect 50308 5958 50338 6010
rect 50362 5958 50372 6010
rect 50372 5958 50418 6010
rect 50442 5958 50488 6010
rect 50488 5958 50498 6010
rect 50522 5958 50552 6010
rect 50552 5958 50578 6010
rect 50282 5956 50338 5958
rect 50362 5956 50418 5958
rect 50442 5956 50498 5958
rect 50522 5956 50578 5958
rect 50282 4922 50338 4924
rect 50362 4922 50418 4924
rect 50442 4922 50498 4924
rect 50522 4922 50578 4924
rect 50282 4870 50308 4922
rect 50308 4870 50338 4922
rect 50362 4870 50372 4922
rect 50372 4870 50418 4922
rect 50442 4870 50488 4922
rect 50488 4870 50498 4922
rect 50522 4870 50552 4922
rect 50552 4870 50578 4922
rect 50282 4868 50338 4870
rect 50362 4868 50418 4870
rect 50442 4868 50498 4870
rect 50522 4868 50578 4870
rect 50282 3834 50338 3836
rect 50362 3834 50418 3836
rect 50442 3834 50498 3836
rect 50522 3834 50578 3836
rect 50282 3782 50308 3834
rect 50308 3782 50338 3834
rect 50362 3782 50372 3834
rect 50372 3782 50418 3834
rect 50442 3782 50488 3834
rect 50488 3782 50498 3834
rect 50522 3782 50552 3834
rect 50552 3782 50578 3834
rect 50282 3780 50338 3782
rect 50362 3780 50418 3782
rect 50442 3780 50498 3782
rect 50522 3780 50578 3782
rect 50282 2746 50338 2748
rect 50362 2746 50418 2748
rect 50442 2746 50498 2748
rect 50522 2746 50578 2748
rect 50282 2694 50308 2746
rect 50308 2694 50338 2746
rect 50362 2694 50372 2746
rect 50372 2694 50418 2746
rect 50442 2694 50488 2746
rect 50488 2694 50498 2746
rect 50522 2694 50552 2746
rect 50552 2694 50578 2746
rect 50282 2692 50338 2694
rect 50362 2692 50418 2694
rect 50442 2692 50498 2694
rect 50522 2692 50578 2694
rect 56764 57976 56820 58032
rect 56948 57976 57004 58032
rect 56396 55800 56452 55856
rect 56856 38800 56912 38856
rect 56764 38664 56820 38720
rect 57132 9560 57188 9616
rect 55660 2896 55716 2952
<< metal3 >>
rect 51239 58034 51305 58037
rect 52251 58034 52317 58037
rect 51239 58032 52317 58034
rect 51239 57976 51244 58032
rect 51300 57976 52256 58032
rect 52312 57976 52317 58032
rect 51239 57974 52317 57976
rect 51239 57971 51305 57974
rect 52251 57971 52317 57974
rect 56759 58034 56825 58037
rect 56943 58034 57009 58037
rect 56759 58032 57009 58034
rect 56759 57976 56764 58032
rect 56820 57976 56948 58032
rect 57004 57976 57009 58032
rect 56759 57974 57009 57976
rect 56759 57971 56825 57974
rect 56943 57971 57009 57974
rect 4190 57696 4510 57697
rect 4190 57632 4198 57696
rect 4262 57632 4278 57696
rect 4342 57632 4358 57696
rect 4422 57632 4438 57696
rect 4502 57632 4510 57696
rect 4190 57631 4510 57632
rect 34910 57696 35230 57697
rect 34910 57632 34918 57696
rect 34982 57632 34998 57696
rect 35062 57632 35078 57696
rect 35142 57632 35158 57696
rect 35222 57632 35230 57696
rect 34910 57631 35230 57632
rect 19550 57152 19870 57153
rect 19550 57088 19558 57152
rect 19622 57088 19638 57152
rect 19702 57088 19718 57152
rect 19782 57088 19798 57152
rect 19862 57088 19870 57152
rect 19550 57087 19870 57088
rect 50270 57152 50590 57153
rect 50270 57088 50278 57152
rect 50342 57088 50358 57152
rect 50422 57088 50438 57152
rect 50502 57088 50518 57152
rect 50582 57088 50590 57152
rect 50270 57087 50590 57088
rect 26951 56810 27017 56813
rect 26724 56808 27017 56810
rect 26724 56752 26956 56808
rect 27012 56752 27017 56808
rect 26724 56750 27017 56752
rect 26724 56674 26784 56750
rect 26951 56747 27017 56750
rect 26859 56674 26925 56677
rect 26724 56672 26925 56674
rect 26724 56616 26864 56672
rect 26920 56616 26925 56672
rect 26724 56614 26925 56616
rect 26859 56611 26925 56614
rect 4190 56608 4510 56609
rect 4190 56544 4198 56608
rect 4262 56544 4278 56608
rect 4342 56544 4358 56608
rect 4422 56544 4438 56608
rect 4502 56544 4510 56608
rect 4190 56543 4510 56544
rect 34910 56608 35230 56609
rect 34910 56544 34918 56608
rect 34982 56544 34998 56608
rect 35062 56544 35078 56608
rect 35142 56544 35158 56608
rect 35222 56544 35230 56608
rect 34910 56543 35230 56544
rect 26675 56402 26741 56405
rect 28147 56402 28213 56405
rect 26675 56400 28213 56402
rect 26675 56344 26680 56400
rect 26736 56344 28152 56400
rect 28208 56344 28213 56400
rect 26675 56342 28213 56344
rect 26675 56339 26741 56342
rect 28147 56339 28213 56342
rect 33759 56402 33825 56405
rect 40199 56402 40265 56405
rect 33759 56400 40265 56402
rect 33759 56344 33764 56400
rect 33820 56344 40204 56400
rect 40260 56344 40265 56400
rect 33759 56342 40265 56344
rect 33759 56339 33825 56342
rect 40199 56339 40265 56342
rect 41119 56402 41185 56405
rect 41487 56402 41553 56405
rect 41119 56400 41553 56402
rect 41119 56344 41124 56400
rect 41180 56344 41492 56400
rect 41548 56344 41553 56400
rect 41119 56342 41553 56344
rect 41119 56339 41185 56342
rect 41487 56339 41553 56342
rect 32471 56266 32537 56269
rect 41303 56266 41369 56269
rect 32471 56264 41369 56266
rect 32471 56208 32476 56264
rect 32532 56208 41308 56264
rect 41364 56208 41369 56264
rect 32471 56206 41369 56208
rect 32471 56203 32537 56206
rect 41303 56203 41369 56206
rect 31643 56130 31709 56133
rect 31827 56130 31893 56133
rect 31643 56128 31893 56130
rect 31643 56072 31648 56128
rect 31704 56072 31832 56128
rect 31888 56072 31893 56128
rect 31643 56070 31893 56072
rect 31643 56067 31709 56070
rect 31827 56067 31893 56070
rect 19550 56064 19870 56065
rect 19550 56000 19558 56064
rect 19622 56000 19638 56064
rect 19702 56000 19718 56064
rect 19782 56000 19798 56064
rect 19862 56000 19870 56064
rect 19550 55999 19870 56000
rect 50270 56064 50590 56065
rect 50270 56000 50278 56064
rect 50342 56000 50358 56064
rect 50422 56000 50438 56064
rect 50502 56000 50518 56064
rect 50582 56000 50590 56064
rect 50270 55999 50590 56000
rect 18487 55858 18553 55861
rect 56391 55858 56457 55861
rect 18487 55856 56457 55858
rect 18487 55800 18492 55856
rect 18548 55800 56396 55856
rect 56452 55800 56457 55856
rect 18487 55798 56457 55800
rect 18487 55795 18553 55798
rect 56391 55795 56457 55798
rect 31551 55722 31617 55725
rect 31735 55722 31801 55725
rect 31551 55720 31801 55722
rect 31551 55664 31556 55720
rect 31612 55664 31740 55720
rect 31796 55664 31801 55720
rect 31551 55662 31801 55664
rect 31551 55659 31617 55662
rect 31735 55659 31801 55662
rect 27411 55586 27477 55589
rect 31183 55586 31249 55589
rect 27411 55584 31249 55586
rect 27411 55528 27416 55584
rect 27472 55528 31188 55584
rect 31244 55528 31249 55584
rect 27411 55526 31249 55528
rect 27411 55523 27477 55526
rect 31183 55523 31249 55526
rect 4190 55520 4510 55521
rect 4190 55456 4198 55520
rect 4262 55456 4278 55520
rect 4342 55456 4358 55520
rect 4422 55456 4438 55520
rect 4502 55456 4510 55520
rect 4190 55455 4510 55456
rect 34910 55520 35230 55521
rect 34910 55456 34918 55520
rect 34982 55456 34998 55520
rect 35062 55456 35078 55520
rect 35142 55456 35158 55520
rect 35222 55456 35230 55520
rect 34910 55455 35230 55456
rect 41303 55450 41369 55453
rect 45443 55450 45509 55453
rect 41303 55448 45509 55450
rect 41303 55392 41308 55448
rect 41364 55392 45448 55448
rect 45504 55392 45509 55448
rect 41303 55390 45509 55392
rect 41303 55387 41369 55390
rect 45443 55387 45509 55390
rect 19550 54976 19870 54977
rect 19550 54912 19558 54976
rect 19622 54912 19638 54976
rect 19702 54912 19718 54976
rect 19782 54912 19798 54976
rect 19862 54912 19870 54976
rect 19550 54911 19870 54912
rect 50270 54976 50590 54977
rect 50270 54912 50278 54976
rect 50342 54912 50358 54976
rect 50422 54912 50438 54976
rect 50502 54912 50518 54976
rect 50582 54912 50590 54976
rect 50270 54911 50590 54912
rect 19315 54634 19381 54637
rect 23547 54634 23613 54637
rect 19315 54632 23613 54634
rect 19315 54576 19320 54632
rect 19376 54576 23552 54632
rect 23608 54576 23613 54632
rect 19315 54574 23613 54576
rect 19315 54571 19381 54574
rect 23547 54571 23613 54574
rect 4190 54432 4510 54433
rect 4190 54368 4198 54432
rect 4262 54368 4278 54432
rect 4342 54368 4358 54432
rect 4422 54368 4438 54432
rect 4502 54368 4510 54432
rect 4190 54367 4510 54368
rect 34910 54432 35230 54433
rect 34910 54368 34918 54432
rect 34982 54368 34998 54432
rect 35062 54368 35078 54432
rect 35142 54368 35158 54432
rect 35222 54368 35230 54432
rect 34910 54367 35230 54368
rect 19550 53888 19870 53889
rect 19550 53824 19558 53888
rect 19622 53824 19638 53888
rect 19702 53824 19718 53888
rect 19782 53824 19798 53888
rect 19862 53824 19870 53888
rect 19550 53823 19870 53824
rect 50270 53888 50590 53889
rect 50270 53824 50278 53888
rect 50342 53824 50358 53888
rect 50422 53824 50438 53888
rect 50502 53824 50518 53888
rect 50582 53824 50590 53888
rect 50270 53823 50590 53824
rect 45535 53818 45601 53821
rect 45719 53818 45785 53821
rect 45535 53816 45785 53818
rect 45535 53760 45540 53816
rect 45596 53760 45724 53816
rect 45780 53760 45785 53816
rect 45535 53758 45785 53760
rect 45535 53755 45601 53758
rect 45719 53755 45785 53758
rect 4190 53344 4510 53345
rect 4190 53280 4198 53344
rect 4262 53280 4278 53344
rect 4342 53280 4358 53344
rect 4422 53280 4438 53344
rect 4502 53280 4510 53344
rect 4190 53279 4510 53280
rect 34910 53344 35230 53345
rect 34910 53280 34918 53344
rect 34982 53280 34998 53344
rect 35062 53280 35078 53344
rect 35142 53280 35158 53344
rect 35222 53280 35230 53344
rect 34910 53279 35230 53280
rect 19550 52800 19870 52801
rect 19550 52736 19558 52800
rect 19622 52736 19638 52800
rect 19702 52736 19718 52800
rect 19782 52736 19798 52800
rect 19862 52736 19870 52800
rect 19550 52735 19870 52736
rect 50270 52800 50590 52801
rect 50270 52736 50278 52800
rect 50342 52736 50358 52800
rect 50422 52736 50438 52800
rect 50502 52736 50518 52800
rect 50582 52736 50590 52800
rect 50270 52735 50590 52736
rect 4190 52256 4510 52257
rect 4190 52192 4198 52256
rect 4262 52192 4278 52256
rect 4342 52192 4358 52256
rect 4422 52192 4438 52256
rect 4502 52192 4510 52256
rect 4190 52191 4510 52192
rect 34910 52256 35230 52257
rect 34910 52192 34918 52256
rect 34982 52192 34998 52256
rect 35062 52192 35078 52256
rect 35142 52192 35158 52256
rect 35222 52192 35230 52256
rect 34910 52191 35230 52192
rect 19550 51712 19870 51713
rect 19550 51648 19558 51712
rect 19622 51648 19638 51712
rect 19702 51648 19718 51712
rect 19782 51648 19798 51712
rect 19862 51648 19870 51712
rect 19550 51647 19870 51648
rect 50270 51712 50590 51713
rect 50270 51648 50278 51712
rect 50342 51648 50358 51712
rect 50422 51648 50438 51712
rect 50502 51648 50518 51712
rect 50582 51648 50590 51712
rect 50270 51647 50590 51648
rect 4190 51168 4510 51169
rect 4190 51104 4198 51168
rect 4262 51104 4278 51168
rect 4342 51104 4358 51168
rect 4422 51104 4438 51168
rect 4502 51104 4510 51168
rect 4190 51103 4510 51104
rect 34910 51168 35230 51169
rect 34910 51104 34918 51168
rect 34982 51104 34998 51168
rect 35062 51104 35078 51168
rect 35142 51104 35158 51168
rect 35222 51104 35230 51168
rect 34910 51103 35230 51104
rect 19550 50624 19870 50625
rect 19550 50560 19558 50624
rect 19622 50560 19638 50624
rect 19702 50560 19718 50624
rect 19782 50560 19798 50624
rect 19862 50560 19870 50624
rect 19550 50559 19870 50560
rect 50270 50624 50590 50625
rect 50270 50560 50278 50624
rect 50342 50560 50358 50624
rect 50422 50560 50438 50624
rect 50502 50560 50518 50624
rect 50582 50560 50590 50624
rect 50270 50559 50590 50560
rect 4190 50080 4510 50081
rect 4190 50016 4198 50080
rect 4262 50016 4278 50080
rect 4342 50016 4358 50080
rect 4422 50016 4438 50080
rect 4502 50016 4510 50080
rect 4190 50015 4510 50016
rect 34910 50080 35230 50081
rect 34910 50016 34918 50080
rect 34982 50016 34998 50080
rect 35062 50016 35078 50080
rect 35142 50016 35158 50080
rect 35222 50016 35230 50080
rect 34910 50015 35230 50016
rect 19550 49536 19870 49537
rect 19550 49472 19558 49536
rect 19622 49472 19638 49536
rect 19702 49472 19718 49536
rect 19782 49472 19798 49536
rect 19862 49472 19870 49536
rect 19550 49471 19870 49472
rect 50270 49536 50590 49537
rect 50270 49472 50278 49536
rect 50342 49472 50358 49536
rect 50422 49472 50438 49536
rect 50502 49472 50518 49536
rect 50582 49472 50590 49536
rect 50270 49471 50590 49472
rect 4190 48992 4510 48993
rect 4190 48928 4198 48992
rect 4262 48928 4278 48992
rect 4342 48928 4358 48992
rect 4422 48928 4438 48992
rect 4502 48928 4510 48992
rect 4190 48927 4510 48928
rect 34910 48992 35230 48993
rect 34910 48928 34918 48992
rect 34982 48928 34998 48992
rect 35062 48928 35078 48992
rect 35142 48928 35158 48992
rect 35222 48928 35230 48992
rect 34910 48927 35230 48928
rect 19550 48448 19870 48449
rect 19550 48384 19558 48448
rect 19622 48384 19638 48448
rect 19702 48384 19718 48448
rect 19782 48384 19798 48448
rect 19862 48384 19870 48448
rect 19550 48383 19870 48384
rect 50270 48448 50590 48449
rect 50270 48384 50278 48448
rect 50342 48384 50358 48448
rect 50422 48384 50438 48448
rect 50502 48384 50518 48448
rect 50582 48384 50590 48448
rect 50270 48383 50590 48384
rect 4190 47904 4510 47905
rect 4190 47840 4198 47904
rect 4262 47840 4278 47904
rect 4342 47840 4358 47904
rect 4422 47840 4438 47904
rect 4502 47840 4510 47904
rect 4190 47839 4510 47840
rect 34910 47904 35230 47905
rect 34910 47840 34918 47904
rect 34982 47840 34998 47904
rect 35062 47840 35078 47904
rect 35142 47840 35158 47904
rect 35222 47840 35230 47904
rect 34910 47839 35230 47840
rect 19550 47360 19870 47361
rect 19550 47296 19558 47360
rect 19622 47296 19638 47360
rect 19702 47296 19718 47360
rect 19782 47296 19798 47360
rect 19862 47296 19870 47360
rect 19550 47295 19870 47296
rect 50270 47360 50590 47361
rect 50270 47296 50278 47360
rect 50342 47296 50358 47360
rect 50422 47296 50438 47360
rect 50502 47296 50518 47360
rect 50582 47296 50590 47360
rect 50270 47295 50590 47296
rect 4190 46816 4510 46817
rect 4190 46752 4198 46816
rect 4262 46752 4278 46816
rect 4342 46752 4358 46816
rect 4422 46752 4438 46816
rect 4502 46752 4510 46816
rect 4190 46751 4510 46752
rect 34910 46816 35230 46817
rect 34910 46752 34918 46816
rect 34982 46752 34998 46816
rect 35062 46752 35078 46816
rect 35142 46752 35158 46816
rect 35222 46752 35230 46816
rect 34910 46751 35230 46752
rect 19550 46272 19870 46273
rect 19550 46208 19558 46272
rect 19622 46208 19638 46272
rect 19702 46208 19718 46272
rect 19782 46208 19798 46272
rect 19862 46208 19870 46272
rect 19550 46207 19870 46208
rect 50270 46272 50590 46273
rect 50270 46208 50278 46272
rect 50342 46208 50358 46272
rect 50422 46208 50438 46272
rect 50502 46208 50518 46272
rect 50582 46208 50590 46272
rect 50270 46207 50590 46208
rect 4190 45728 4510 45729
rect 4190 45664 4198 45728
rect 4262 45664 4278 45728
rect 4342 45664 4358 45728
rect 4422 45664 4438 45728
rect 4502 45664 4510 45728
rect 4190 45663 4510 45664
rect 34910 45728 35230 45729
rect 34910 45664 34918 45728
rect 34982 45664 34998 45728
rect 35062 45664 35078 45728
rect 35142 45664 35158 45728
rect 35222 45664 35230 45728
rect 34910 45663 35230 45664
rect 19550 45184 19870 45185
rect 19550 45120 19558 45184
rect 19622 45120 19638 45184
rect 19702 45120 19718 45184
rect 19782 45120 19798 45184
rect 19862 45120 19870 45184
rect 19550 45119 19870 45120
rect 50270 45184 50590 45185
rect 50270 45120 50278 45184
rect 50342 45120 50358 45184
rect 50422 45120 50438 45184
rect 50502 45120 50518 45184
rect 50582 45120 50590 45184
rect 50270 45119 50590 45120
rect 4190 44640 4510 44641
rect 4190 44576 4198 44640
rect 4262 44576 4278 44640
rect 4342 44576 4358 44640
rect 4422 44576 4438 44640
rect 4502 44576 4510 44640
rect 4190 44575 4510 44576
rect 34910 44640 35230 44641
rect 34910 44576 34918 44640
rect 34982 44576 34998 44640
rect 35062 44576 35078 44640
rect 35142 44576 35158 44640
rect 35222 44576 35230 44640
rect 34910 44575 35230 44576
rect 22995 44162 23061 44165
rect 23179 44162 23245 44165
rect 38819 44164 38885 44165
rect 38819 44162 38866 44164
rect 22995 44160 23245 44162
rect 22995 44104 23000 44160
rect 23056 44104 23184 44160
rect 23240 44104 23245 44160
rect 22995 44102 23245 44104
rect 38774 44160 38866 44162
rect 38774 44104 38824 44160
rect 38774 44102 38866 44104
rect 22995 44099 23061 44102
rect 23179 44099 23245 44102
rect 38819 44100 38866 44102
rect 38930 44100 38936 44164
rect 38819 44099 38885 44100
rect 19550 44096 19870 44097
rect 19550 44032 19558 44096
rect 19622 44032 19638 44096
rect 19702 44032 19718 44096
rect 19782 44032 19798 44096
rect 19862 44032 19870 44096
rect 19550 44031 19870 44032
rect 50270 44096 50590 44097
rect 50270 44032 50278 44096
rect 50342 44032 50358 44096
rect 50422 44032 50438 44096
rect 50502 44032 50518 44096
rect 50582 44032 50590 44096
rect 50270 44031 50590 44032
rect 4190 43552 4510 43553
rect 4190 43488 4198 43552
rect 4262 43488 4278 43552
rect 4342 43488 4358 43552
rect 4422 43488 4438 43552
rect 4502 43488 4510 43552
rect 4190 43487 4510 43488
rect 34910 43552 35230 43553
rect 34910 43488 34918 43552
rect 34982 43488 34998 43552
rect 35062 43488 35078 43552
rect 35142 43488 35158 43552
rect 35222 43488 35230 43552
rect 34910 43487 35230 43488
rect 19550 43008 19870 43009
rect 19550 42944 19558 43008
rect 19622 42944 19638 43008
rect 19702 42944 19718 43008
rect 19782 42944 19798 43008
rect 19862 42944 19870 43008
rect 19550 42943 19870 42944
rect 50270 43008 50590 43009
rect 50270 42944 50278 43008
rect 50342 42944 50358 43008
rect 50422 42944 50438 43008
rect 50502 42944 50518 43008
rect 50582 42944 50590 43008
rect 50270 42943 50590 42944
rect 4190 42464 4510 42465
rect 4190 42400 4198 42464
rect 4262 42400 4278 42464
rect 4342 42400 4358 42464
rect 4422 42400 4438 42464
rect 4502 42400 4510 42464
rect 4190 42399 4510 42400
rect 34910 42464 35230 42465
rect 34910 42400 34918 42464
rect 34982 42400 34998 42464
rect 35062 42400 35078 42464
rect 35142 42400 35158 42464
rect 35222 42400 35230 42464
rect 34910 42399 35230 42400
rect 19550 41920 19870 41921
rect 19550 41856 19558 41920
rect 19622 41856 19638 41920
rect 19702 41856 19718 41920
rect 19782 41856 19798 41920
rect 19862 41856 19870 41920
rect 19550 41855 19870 41856
rect 50270 41920 50590 41921
rect 50270 41856 50278 41920
rect 50342 41856 50358 41920
rect 50422 41856 50438 41920
rect 50502 41856 50518 41920
rect 50582 41856 50590 41920
rect 50270 41855 50590 41856
rect 4190 41376 4510 41377
rect 4190 41312 4198 41376
rect 4262 41312 4278 41376
rect 4342 41312 4358 41376
rect 4422 41312 4438 41376
rect 4502 41312 4510 41376
rect 4190 41311 4510 41312
rect 34910 41376 35230 41377
rect 34910 41312 34918 41376
rect 34982 41312 34998 41376
rect 35062 41312 35078 41376
rect 35142 41312 35158 41376
rect 35222 41312 35230 41376
rect 34910 41311 35230 41312
rect 19550 40832 19870 40833
rect 19550 40768 19558 40832
rect 19622 40768 19638 40832
rect 19702 40768 19718 40832
rect 19782 40768 19798 40832
rect 19862 40768 19870 40832
rect 19550 40767 19870 40768
rect 50270 40832 50590 40833
rect 50270 40768 50278 40832
rect 50342 40768 50358 40832
rect 50422 40768 50438 40832
rect 50502 40768 50518 40832
rect 50582 40768 50590 40832
rect 50270 40767 50590 40768
rect 4190 40288 4510 40289
rect 4190 40224 4198 40288
rect 4262 40224 4278 40288
rect 4342 40224 4358 40288
rect 4422 40224 4438 40288
rect 4502 40224 4510 40288
rect 4190 40223 4510 40224
rect 34910 40288 35230 40289
rect 34910 40224 34918 40288
rect 34982 40224 34998 40288
rect 35062 40224 35078 40288
rect 35142 40224 35158 40288
rect 35222 40224 35230 40288
rect 34910 40223 35230 40224
rect 19550 39744 19870 39745
rect 19550 39680 19558 39744
rect 19622 39680 19638 39744
rect 19702 39680 19718 39744
rect 19782 39680 19798 39744
rect 19862 39680 19870 39744
rect 19550 39679 19870 39680
rect 50270 39744 50590 39745
rect 50270 39680 50278 39744
rect 50342 39680 50358 39744
rect 50422 39680 50438 39744
rect 50502 39680 50518 39744
rect 50582 39680 50590 39744
rect 50270 39679 50590 39680
rect 4190 39200 4510 39201
rect 4190 39136 4198 39200
rect 4262 39136 4278 39200
rect 4342 39136 4358 39200
rect 4422 39136 4438 39200
rect 4502 39136 4510 39200
rect 4190 39135 4510 39136
rect 34910 39200 35230 39201
rect 34910 39136 34918 39200
rect 34982 39136 34998 39200
rect 35062 39136 35078 39200
rect 35142 39136 35158 39200
rect 35222 39136 35230 39200
rect 34910 39135 35230 39136
rect 56851 38858 56917 38861
rect 56716 38856 56917 38858
rect 56716 38800 56856 38856
rect 56912 38800 56917 38856
rect 56716 38798 56917 38800
rect 56716 38725 56776 38798
rect 56851 38795 56917 38798
rect 24099 38722 24165 38725
rect 29343 38722 29409 38725
rect 24099 38720 24208 38722
rect 24099 38664 24104 38720
rect 24160 38664 24208 38720
rect 24099 38659 24208 38664
rect 19550 38656 19870 38657
rect 19550 38592 19558 38656
rect 19622 38592 19638 38656
rect 19702 38592 19718 38656
rect 19782 38592 19798 38656
rect 19862 38592 19870 38656
rect 19550 38591 19870 38592
rect 24148 38589 24208 38659
rect 24099 38584 24208 38589
rect 24099 38528 24104 38584
rect 24160 38528 24208 38584
rect 24099 38526 24208 38528
rect 29116 38720 29409 38722
rect 29116 38664 29348 38720
rect 29404 38664 29409 38720
rect 29116 38662 29409 38664
rect 56716 38720 56825 38725
rect 56716 38664 56764 38720
rect 56820 38664 56825 38720
rect 56716 38662 56825 38664
rect 29116 38586 29176 38662
rect 29343 38659 29409 38662
rect 56759 38659 56825 38662
rect 50270 38656 50590 38657
rect 50270 38592 50278 38656
rect 50342 38592 50358 38656
rect 50422 38592 50438 38656
rect 50502 38592 50518 38656
rect 50582 38592 50590 38656
rect 50270 38591 50590 38592
rect 29251 38586 29317 38589
rect 29116 38584 29317 38586
rect 29116 38528 29256 38584
rect 29312 38528 29317 38584
rect 29116 38526 29317 38528
rect 24099 38523 24165 38526
rect 29251 38523 29317 38526
rect 4190 38112 4510 38113
rect 4190 38048 4198 38112
rect 4262 38048 4278 38112
rect 4342 38048 4358 38112
rect 4422 38048 4438 38112
rect 4502 38048 4510 38112
rect 4190 38047 4510 38048
rect 34910 38112 35230 38113
rect 34910 38048 34918 38112
rect 34982 38048 34998 38112
rect 35062 38048 35078 38112
rect 35142 38048 35158 38112
rect 35222 38048 35230 38112
rect 34910 38047 35230 38048
rect 19550 37568 19870 37569
rect 19550 37504 19558 37568
rect 19622 37504 19638 37568
rect 19702 37504 19718 37568
rect 19782 37504 19798 37568
rect 19862 37504 19870 37568
rect 19550 37503 19870 37504
rect 50270 37568 50590 37569
rect 50270 37504 50278 37568
rect 50342 37504 50358 37568
rect 50422 37504 50438 37568
rect 50502 37504 50518 37568
rect 50582 37504 50590 37568
rect 50270 37503 50590 37504
rect 4190 37024 4510 37025
rect 4190 36960 4198 37024
rect 4262 36960 4278 37024
rect 4342 36960 4358 37024
rect 4422 36960 4438 37024
rect 4502 36960 4510 37024
rect 4190 36959 4510 36960
rect 34910 37024 35230 37025
rect 34910 36960 34918 37024
rect 34982 36960 34998 37024
rect 35062 36960 35078 37024
rect 35142 36960 35158 37024
rect 35222 36960 35230 37024
rect 34910 36959 35230 36960
rect 19550 36480 19870 36481
rect 19550 36416 19558 36480
rect 19622 36416 19638 36480
rect 19702 36416 19718 36480
rect 19782 36416 19798 36480
rect 19862 36416 19870 36480
rect 19550 36415 19870 36416
rect 50270 36480 50590 36481
rect 50270 36416 50278 36480
rect 50342 36416 50358 36480
rect 50422 36416 50438 36480
rect 50502 36416 50518 36480
rect 50582 36416 50590 36480
rect 50270 36415 50590 36416
rect 4190 35936 4510 35937
rect 4190 35872 4198 35936
rect 4262 35872 4278 35936
rect 4342 35872 4358 35936
rect 4422 35872 4438 35936
rect 4502 35872 4510 35936
rect 4190 35871 4510 35872
rect 34910 35936 35230 35937
rect 34910 35872 34918 35936
rect 34982 35872 34998 35936
rect 35062 35872 35078 35936
rect 35142 35872 35158 35936
rect 35222 35872 35230 35936
rect 34910 35871 35230 35872
rect 19550 35392 19870 35393
rect 19550 35328 19558 35392
rect 19622 35328 19638 35392
rect 19702 35328 19718 35392
rect 19782 35328 19798 35392
rect 19862 35328 19870 35392
rect 19550 35327 19870 35328
rect 50270 35392 50590 35393
rect 50270 35328 50278 35392
rect 50342 35328 50358 35392
rect 50422 35328 50438 35392
rect 50502 35328 50518 35392
rect 50582 35328 50590 35392
rect 50270 35327 50590 35328
rect 4190 34848 4510 34849
rect 4190 34784 4198 34848
rect 4262 34784 4278 34848
rect 4342 34784 4358 34848
rect 4422 34784 4438 34848
rect 4502 34784 4510 34848
rect 4190 34783 4510 34784
rect 34910 34848 35230 34849
rect 34910 34784 34918 34848
rect 34982 34784 34998 34848
rect 35062 34784 35078 34848
rect 35142 34784 35158 34848
rect 35222 34784 35230 34848
rect 34910 34783 35230 34784
rect 45535 34506 45601 34509
rect 45719 34506 45785 34509
rect 45535 34504 45785 34506
rect 45535 34448 45540 34504
rect 45596 34448 45724 34504
rect 45780 34448 45785 34504
rect 45535 34446 45785 34448
rect 45535 34443 45601 34446
rect 45719 34443 45785 34446
rect 19550 34304 19870 34305
rect 19550 34240 19558 34304
rect 19622 34240 19638 34304
rect 19702 34240 19718 34304
rect 19782 34240 19798 34304
rect 19862 34240 19870 34304
rect 19550 34239 19870 34240
rect 50270 34304 50590 34305
rect 50270 34240 50278 34304
rect 50342 34240 50358 34304
rect 50422 34240 50438 34304
rect 50502 34240 50518 34304
rect 50582 34240 50590 34304
rect 50270 34239 50590 34240
rect 4190 33760 4510 33761
rect 4190 33696 4198 33760
rect 4262 33696 4278 33760
rect 4342 33696 4358 33760
rect 4422 33696 4438 33760
rect 4502 33696 4510 33760
rect 4190 33695 4510 33696
rect 34910 33760 35230 33761
rect 34910 33696 34918 33760
rect 34982 33696 34998 33760
rect 35062 33696 35078 33760
rect 35142 33696 35158 33760
rect 35222 33696 35230 33760
rect 34910 33695 35230 33696
rect 19550 33216 19870 33217
rect 19550 33152 19558 33216
rect 19622 33152 19638 33216
rect 19702 33152 19718 33216
rect 19782 33152 19798 33216
rect 19862 33152 19870 33216
rect 19550 33151 19870 33152
rect 50270 33216 50590 33217
rect 50270 33152 50278 33216
rect 50342 33152 50358 33216
rect 50422 33152 50438 33216
rect 50502 33152 50518 33216
rect 50582 33152 50590 33216
rect 50270 33151 50590 33152
rect 4190 32672 4510 32673
rect 4190 32608 4198 32672
rect 4262 32608 4278 32672
rect 4342 32608 4358 32672
rect 4422 32608 4438 32672
rect 4502 32608 4510 32672
rect 4190 32607 4510 32608
rect 34910 32672 35230 32673
rect 34910 32608 34918 32672
rect 34982 32608 34998 32672
rect 35062 32608 35078 32672
rect 35142 32608 35158 32672
rect 35222 32608 35230 32672
rect 34910 32607 35230 32608
rect 19550 32128 19870 32129
rect 19550 32064 19558 32128
rect 19622 32064 19638 32128
rect 19702 32064 19718 32128
rect 19782 32064 19798 32128
rect 19862 32064 19870 32128
rect 19550 32063 19870 32064
rect 50270 32128 50590 32129
rect 50270 32064 50278 32128
rect 50342 32064 50358 32128
rect 50422 32064 50438 32128
rect 50502 32064 50518 32128
rect 50582 32064 50590 32128
rect 50270 32063 50590 32064
rect 4190 31584 4510 31585
rect 4190 31520 4198 31584
rect 4262 31520 4278 31584
rect 4342 31520 4358 31584
rect 4422 31520 4438 31584
rect 4502 31520 4510 31584
rect 4190 31519 4510 31520
rect 34910 31584 35230 31585
rect 34910 31520 34918 31584
rect 34982 31520 34998 31584
rect 35062 31520 35078 31584
rect 35142 31520 35158 31584
rect 35222 31520 35230 31584
rect 34910 31519 35230 31520
rect 19550 31040 19870 31041
rect 19550 30976 19558 31040
rect 19622 30976 19638 31040
rect 19702 30976 19718 31040
rect 19782 30976 19798 31040
rect 19862 30976 19870 31040
rect 19550 30975 19870 30976
rect 50270 31040 50590 31041
rect 50270 30976 50278 31040
rect 50342 30976 50358 31040
rect 50422 30976 50438 31040
rect 50502 30976 50518 31040
rect 50582 30976 50590 31040
rect 50270 30975 50590 30976
rect 4190 30496 4510 30497
rect 4190 30432 4198 30496
rect 4262 30432 4278 30496
rect 4342 30432 4358 30496
rect 4422 30432 4438 30496
rect 4502 30432 4510 30496
rect 4190 30431 4510 30432
rect 34910 30496 35230 30497
rect 34910 30432 34918 30496
rect 34982 30432 34998 30496
rect 35062 30432 35078 30496
rect 35142 30432 35158 30496
rect 35222 30432 35230 30496
rect 34910 30431 35230 30432
rect 19550 29952 19870 29953
rect 19550 29888 19558 29952
rect 19622 29888 19638 29952
rect 19702 29888 19718 29952
rect 19782 29888 19798 29952
rect 19862 29888 19870 29952
rect 19550 29887 19870 29888
rect 50270 29952 50590 29953
rect 50270 29888 50278 29952
rect 50342 29888 50358 29952
rect 50422 29888 50438 29952
rect 50502 29888 50518 29952
rect 50582 29888 50590 29952
rect 50270 29887 50590 29888
rect 4190 29408 4510 29409
rect 4190 29344 4198 29408
rect 4262 29344 4278 29408
rect 4342 29344 4358 29408
rect 4422 29344 4438 29408
rect 4502 29344 4510 29408
rect 4190 29343 4510 29344
rect 34910 29408 35230 29409
rect 34910 29344 34918 29408
rect 34982 29344 34998 29408
rect 35062 29344 35078 29408
rect 35142 29344 35158 29408
rect 35222 29344 35230 29408
rect 34910 29343 35230 29344
rect 18855 29066 18921 29069
rect 18812 29064 18921 29066
rect 18812 29008 18860 29064
rect 18916 29008 18921 29064
rect 18812 29003 18921 29008
rect 18812 28930 18872 29003
rect 18947 28930 19013 28933
rect 18812 28928 19013 28930
rect 18812 28872 18952 28928
rect 19008 28872 19013 28928
rect 18812 28870 19013 28872
rect 18947 28867 19013 28870
rect 19550 28864 19870 28865
rect 19550 28800 19558 28864
rect 19622 28800 19638 28864
rect 19702 28800 19718 28864
rect 19782 28800 19798 28864
rect 19862 28800 19870 28864
rect 19550 28799 19870 28800
rect 50270 28864 50590 28865
rect 50270 28800 50278 28864
rect 50342 28800 50358 28864
rect 50422 28800 50438 28864
rect 50502 28800 50518 28864
rect 50582 28800 50590 28864
rect 50270 28799 50590 28800
rect 4190 28320 4510 28321
rect 4190 28256 4198 28320
rect 4262 28256 4278 28320
rect 4342 28256 4358 28320
rect 4422 28256 4438 28320
rect 4502 28256 4510 28320
rect 4190 28255 4510 28256
rect 34910 28320 35230 28321
rect 34910 28256 34918 28320
rect 34982 28256 34998 28320
rect 35062 28256 35078 28320
rect 35142 28256 35158 28320
rect 35222 28256 35230 28320
rect 34910 28255 35230 28256
rect 19550 27776 19870 27777
rect 19550 27712 19558 27776
rect 19622 27712 19638 27776
rect 19702 27712 19718 27776
rect 19782 27712 19798 27776
rect 19862 27712 19870 27776
rect 19550 27711 19870 27712
rect 50270 27776 50590 27777
rect 50270 27712 50278 27776
rect 50342 27712 50358 27776
rect 50422 27712 50438 27776
rect 50502 27712 50518 27776
rect 50582 27712 50590 27776
rect 50270 27711 50590 27712
rect 4190 27232 4510 27233
rect 4190 27168 4198 27232
rect 4262 27168 4278 27232
rect 4342 27168 4358 27232
rect 4422 27168 4438 27232
rect 4502 27168 4510 27232
rect 4190 27167 4510 27168
rect 34910 27232 35230 27233
rect 34910 27168 34918 27232
rect 34982 27168 34998 27232
rect 35062 27168 35078 27232
rect 35142 27168 35158 27232
rect 35222 27168 35230 27232
rect 34910 27167 35230 27168
rect 19550 26688 19870 26689
rect 19550 26624 19558 26688
rect 19622 26624 19638 26688
rect 19702 26624 19718 26688
rect 19782 26624 19798 26688
rect 19862 26624 19870 26688
rect 19550 26623 19870 26624
rect 50270 26688 50590 26689
rect 50270 26624 50278 26688
rect 50342 26624 50358 26688
rect 50422 26624 50438 26688
rect 50502 26624 50518 26688
rect 50582 26624 50590 26688
rect 50270 26623 50590 26624
rect 38860 26284 38866 26348
rect 38930 26346 38936 26348
rect 39003 26346 39069 26349
rect 38930 26344 39069 26346
rect 38930 26288 39008 26344
rect 39064 26288 39069 26344
rect 38930 26286 39069 26288
rect 38930 26284 38936 26286
rect 39003 26283 39069 26286
rect 4190 26144 4510 26145
rect 4190 26080 4198 26144
rect 4262 26080 4278 26144
rect 4342 26080 4358 26144
rect 4422 26080 4438 26144
rect 4502 26080 4510 26144
rect 4190 26079 4510 26080
rect 34910 26144 35230 26145
rect 34910 26080 34918 26144
rect 34982 26080 34998 26144
rect 35062 26080 35078 26144
rect 35142 26080 35158 26144
rect 35222 26080 35230 26144
rect 34910 26079 35230 26080
rect 19550 25600 19870 25601
rect 19550 25536 19558 25600
rect 19622 25536 19638 25600
rect 19702 25536 19718 25600
rect 19782 25536 19798 25600
rect 19862 25536 19870 25600
rect 19550 25535 19870 25536
rect 50270 25600 50590 25601
rect 50270 25536 50278 25600
rect 50342 25536 50358 25600
rect 50422 25536 50438 25600
rect 50502 25536 50518 25600
rect 50582 25536 50590 25600
rect 50270 25535 50590 25536
rect 4190 25056 4510 25057
rect 4190 24992 4198 25056
rect 4262 24992 4278 25056
rect 4342 24992 4358 25056
rect 4422 24992 4438 25056
rect 4502 24992 4510 25056
rect 4190 24991 4510 24992
rect 34910 25056 35230 25057
rect 34910 24992 34918 25056
rect 34982 24992 34998 25056
rect 35062 24992 35078 25056
rect 35142 24992 35158 25056
rect 35222 24992 35230 25056
rect 34910 24991 35230 24992
rect 45351 24850 45417 24853
rect 45719 24850 45785 24853
rect 45351 24848 45785 24850
rect 45351 24792 45356 24848
rect 45412 24792 45724 24848
rect 45780 24792 45785 24848
rect 45351 24790 45785 24792
rect 45351 24787 45417 24790
rect 45719 24787 45785 24790
rect 19550 24512 19870 24513
rect 19550 24448 19558 24512
rect 19622 24448 19638 24512
rect 19702 24448 19718 24512
rect 19782 24448 19798 24512
rect 19862 24448 19870 24512
rect 19550 24447 19870 24448
rect 50270 24512 50590 24513
rect 50270 24448 50278 24512
rect 50342 24448 50358 24512
rect 50422 24448 50438 24512
rect 50502 24448 50518 24512
rect 50582 24448 50590 24512
rect 50270 24447 50590 24448
rect 4190 23968 4510 23969
rect 4190 23904 4198 23968
rect 4262 23904 4278 23968
rect 4342 23904 4358 23968
rect 4422 23904 4438 23968
rect 4502 23904 4510 23968
rect 4190 23903 4510 23904
rect 34910 23968 35230 23969
rect 34910 23904 34918 23968
rect 34982 23904 34998 23968
rect 35062 23904 35078 23968
rect 35142 23904 35158 23968
rect 35222 23904 35230 23968
rect 34910 23903 35230 23904
rect 19550 23424 19870 23425
rect 19550 23360 19558 23424
rect 19622 23360 19638 23424
rect 19702 23360 19718 23424
rect 19782 23360 19798 23424
rect 19862 23360 19870 23424
rect 19550 23359 19870 23360
rect 50270 23424 50590 23425
rect 50270 23360 50278 23424
rect 50342 23360 50358 23424
rect 50422 23360 50438 23424
rect 50502 23360 50518 23424
rect 50582 23360 50590 23424
rect 50270 23359 50590 23360
rect 23404 23292 23410 23356
rect 23474 23354 23480 23356
rect 23547 23354 23613 23357
rect 23474 23352 23613 23354
rect 23474 23296 23552 23352
rect 23608 23296 23613 23352
rect 23474 23294 23613 23296
rect 23474 23292 23480 23294
rect 23547 23291 23613 23294
rect 4190 22880 4510 22881
rect 4190 22816 4198 22880
rect 4262 22816 4278 22880
rect 4342 22816 4358 22880
rect 4422 22816 4438 22880
rect 4502 22816 4510 22880
rect 4190 22815 4510 22816
rect 34910 22880 35230 22881
rect 34910 22816 34918 22880
rect 34982 22816 34998 22880
rect 35062 22816 35078 22880
rect 35142 22816 35158 22880
rect 35222 22816 35230 22880
rect 34910 22815 35230 22816
rect 19550 22336 19870 22337
rect 19550 22272 19558 22336
rect 19622 22272 19638 22336
rect 19702 22272 19718 22336
rect 19782 22272 19798 22336
rect 19862 22272 19870 22336
rect 19550 22271 19870 22272
rect 50270 22336 50590 22337
rect 50270 22272 50278 22336
rect 50342 22272 50358 22336
rect 50422 22272 50438 22336
rect 50502 22272 50518 22336
rect 50582 22272 50590 22336
rect 50270 22271 50590 22272
rect 4190 21792 4510 21793
rect 4190 21728 4198 21792
rect 4262 21728 4278 21792
rect 4342 21728 4358 21792
rect 4422 21728 4438 21792
rect 4502 21728 4510 21792
rect 4190 21727 4510 21728
rect 34910 21792 35230 21793
rect 34910 21728 34918 21792
rect 34982 21728 34998 21792
rect 35062 21728 35078 21792
rect 35142 21728 35158 21792
rect 35222 21728 35230 21792
rect 34910 21727 35230 21728
rect 19550 21248 19870 21249
rect 19550 21184 19558 21248
rect 19622 21184 19638 21248
rect 19702 21184 19718 21248
rect 19782 21184 19798 21248
rect 19862 21184 19870 21248
rect 19550 21183 19870 21184
rect 50270 21248 50590 21249
rect 50270 21184 50278 21248
rect 50342 21184 50358 21248
rect 50422 21184 50438 21248
rect 50502 21184 50518 21248
rect 50582 21184 50590 21248
rect 50270 21183 50590 21184
rect 4190 20704 4510 20705
rect 4190 20640 4198 20704
rect 4262 20640 4278 20704
rect 4342 20640 4358 20704
rect 4422 20640 4438 20704
rect 4502 20640 4510 20704
rect 4190 20639 4510 20640
rect 34910 20704 35230 20705
rect 34910 20640 34918 20704
rect 34982 20640 34998 20704
rect 35062 20640 35078 20704
rect 35142 20640 35158 20704
rect 35222 20640 35230 20704
rect 34910 20639 35230 20640
rect 19550 20160 19870 20161
rect 19550 20096 19558 20160
rect 19622 20096 19638 20160
rect 19702 20096 19718 20160
rect 19782 20096 19798 20160
rect 19862 20096 19870 20160
rect 19550 20095 19870 20096
rect 50270 20160 50590 20161
rect 50270 20096 50278 20160
rect 50342 20096 50358 20160
rect 50422 20096 50438 20160
rect 50502 20096 50518 20160
rect 50582 20096 50590 20160
rect 50270 20095 50590 20096
rect 4190 19616 4510 19617
rect 4190 19552 4198 19616
rect 4262 19552 4278 19616
rect 4342 19552 4358 19616
rect 4422 19552 4438 19616
rect 4502 19552 4510 19616
rect 4190 19551 4510 19552
rect 34910 19616 35230 19617
rect 34910 19552 34918 19616
rect 34982 19552 34998 19616
rect 35062 19552 35078 19616
rect 35142 19552 35158 19616
rect 35222 19552 35230 19616
rect 34910 19551 35230 19552
rect 8459 19410 8525 19413
rect 15543 19410 15609 19413
rect 8459 19408 15609 19410
rect 8459 19352 8464 19408
rect 8520 19352 15548 19408
rect 15604 19352 15609 19408
rect 8459 19350 15609 19352
rect 8459 19347 8525 19350
rect 15543 19347 15609 19350
rect 48295 19274 48361 19277
rect 48295 19272 48496 19274
rect 48295 19216 48300 19272
rect 48356 19216 48496 19272
rect 48295 19214 48496 19216
rect 48295 19211 48361 19214
rect 48436 19141 48496 19214
rect 8183 19138 8249 19141
rect 8919 19138 8985 19141
rect 8183 19136 8985 19138
rect 8183 19080 8188 19136
rect 8244 19080 8924 19136
rect 8980 19080 8985 19136
rect 8183 19078 8985 19080
rect 8183 19075 8249 19078
rect 8919 19075 8985 19078
rect 48387 19136 48496 19141
rect 48387 19080 48392 19136
rect 48448 19080 48496 19136
rect 48387 19078 48496 19080
rect 48387 19075 48453 19078
rect 19550 19072 19870 19073
rect 19550 19008 19558 19072
rect 19622 19008 19638 19072
rect 19702 19008 19718 19072
rect 19782 19008 19798 19072
rect 19862 19008 19870 19072
rect 19550 19007 19870 19008
rect 50270 19072 50590 19073
rect 50270 19008 50278 19072
rect 50342 19008 50358 19072
rect 50422 19008 50438 19072
rect 50502 19008 50518 19072
rect 50582 19008 50590 19072
rect 50270 19007 50590 19008
rect 4190 18528 4510 18529
rect 4190 18464 4198 18528
rect 4262 18464 4278 18528
rect 4342 18464 4358 18528
rect 4422 18464 4438 18528
rect 4502 18464 4510 18528
rect 4190 18463 4510 18464
rect 34910 18528 35230 18529
rect 34910 18464 34918 18528
rect 34982 18464 34998 18528
rect 35062 18464 35078 18528
rect 35142 18464 35158 18528
rect 35222 18464 35230 18528
rect 34910 18463 35230 18464
rect 18855 18050 18921 18053
rect 18855 18048 19056 18050
rect 18855 17992 18860 18048
rect 18916 17992 19056 18048
rect 18855 17990 19056 17992
rect 18855 17987 18921 17990
rect 18996 17917 19056 17990
rect 19550 17984 19870 17985
rect 19550 17920 19558 17984
rect 19622 17920 19638 17984
rect 19702 17920 19718 17984
rect 19782 17920 19798 17984
rect 19862 17920 19870 17984
rect 19550 17919 19870 17920
rect 50270 17984 50590 17985
rect 50270 17920 50278 17984
rect 50342 17920 50358 17984
rect 50422 17920 50438 17984
rect 50502 17920 50518 17984
rect 50582 17920 50590 17984
rect 50270 17919 50590 17920
rect 18947 17912 19056 17917
rect 18947 17856 18952 17912
rect 19008 17856 19056 17912
rect 18947 17854 19056 17856
rect 18947 17851 19013 17854
rect 19315 17506 19381 17509
rect 24559 17506 24625 17509
rect 19315 17504 24625 17506
rect 19315 17448 19320 17504
rect 19376 17448 24564 17504
rect 24620 17448 24625 17504
rect 19315 17446 24625 17448
rect 19315 17443 19381 17446
rect 24559 17443 24625 17446
rect 4190 17440 4510 17441
rect 4190 17376 4198 17440
rect 4262 17376 4278 17440
rect 4342 17376 4358 17440
rect 4422 17376 4438 17440
rect 4502 17376 4510 17440
rect 4190 17375 4510 17376
rect 34910 17440 35230 17441
rect 34910 17376 34918 17440
rect 34982 17376 34998 17440
rect 35062 17376 35078 17440
rect 35142 17376 35158 17440
rect 35222 17376 35230 17440
rect 34910 17375 35230 17376
rect 9195 17234 9261 17237
rect 23363 17234 23429 17237
rect 9195 17232 23429 17234
rect 9195 17176 9200 17232
rect 9256 17176 23368 17232
rect 23424 17176 23429 17232
rect 9195 17174 23429 17176
rect 9195 17171 9261 17174
rect 23363 17171 23429 17174
rect 19550 16896 19870 16897
rect 19550 16832 19558 16896
rect 19622 16832 19638 16896
rect 19702 16832 19718 16896
rect 19782 16832 19798 16896
rect 19862 16832 19870 16896
rect 19550 16831 19870 16832
rect 50270 16896 50590 16897
rect 50270 16832 50278 16896
rect 50342 16832 50358 16896
rect 50422 16832 50438 16896
rect 50502 16832 50518 16896
rect 50582 16832 50590 16896
rect 50270 16831 50590 16832
rect 38727 16690 38793 16693
rect 38727 16688 38928 16690
rect 38727 16632 38732 16688
rect 38788 16632 38928 16688
rect 38727 16630 38928 16632
rect 38727 16627 38793 16630
rect 37347 16554 37413 16557
rect 38868 16554 38928 16630
rect 37347 16552 38928 16554
rect 37347 16496 37352 16552
rect 37408 16496 38928 16552
rect 37347 16494 38928 16496
rect 37347 16491 37413 16494
rect 4190 16352 4510 16353
rect 4190 16288 4198 16352
rect 4262 16288 4278 16352
rect 4342 16288 4358 16352
rect 4422 16288 4438 16352
rect 4502 16288 4510 16352
rect 4190 16287 4510 16288
rect 34910 16352 35230 16353
rect 34910 16288 34918 16352
rect 34982 16288 34998 16352
rect 35062 16288 35078 16352
rect 35142 16288 35158 16352
rect 35222 16288 35230 16352
rect 34910 16287 35230 16288
rect 15316 15950 20160 16010
rect 15175 15874 15241 15877
rect 15316 15874 15376 15950
rect 15175 15872 15376 15874
rect 15175 15816 15180 15872
rect 15236 15816 15376 15872
rect 15175 15814 15376 15816
rect 20100 15874 20160 15950
rect 24743 15874 24809 15877
rect 20100 15872 24809 15874
rect 20100 15816 24748 15872
rect 24804 15816 24809 15872
rect 20100 15814 24809 15816
rect 15175 15811 15241 15814
rect 24743 15811 24809 15814
rect 19550 15808 19870 15809
rect 19550 15744 19558 15808
rect 19622 15744 19638 15808
rect 19702 15744 19718 15808
rect 19782 15744 19798 15808
rect 19862 15744 19870 15808
rect 19550 15743 19870 15744
rect 50270 15808 50590 15809
rect 50270 15744 50278 15808
rect 50342 15744 50358 15808
rect 50422 15744 50438 15808
rect 50502 15744 50518 15808
rect 50582 15744 50590 15808
rect 50270 15743 50590 15744
rect 4190 15264 4510 15265
rect 4190 15200 4198 15264
rect 4262 15200 4278 15264
rect 4342 15200 4358 15264
rect 4422 15200 4438 15264
rect 4502 15200 4510 15264
rect 4190 15199 4510 15200
rect 34910 15264 35230 15265
rect 34910 15200 34918 15264
rect 34982 15200 34998 15264
rect 35062 15200 35078 15264
rect 35142 15200 35158 15264
rect 35222 15200 35230 15264
rect 34910 15199 35230 15200
rect 23271 15194 23337 15197
rect 23404 15194 23410 15196
rect 23271 15192 23410 15194
rect 23271 15136 23276 15192
rect 23332 15136 23410 15192
rect 23271 15134 23410 15136
rect 23271 15131 23337 15134
rect 23404 15132 23410 15134
rect 23474 15132 23480 15196
rect 19550 14720 19870 14721
rect 19550 14656 19558 14720
rect 19622 14656 19638 14720
rect 19702 14656 19718 14720
rect 19782 14656 19798 14720
rect 19862 14656 19870 14720
rect 19550 14655 19870 14656
rect 50270 14720 50590 14721
rect 50270 14656 50278 14720
rect 50342 14656 50358 14720
rect 50422 14656 50438 14720
rect 50502 14656 50518 14720
rect 50582 14656 50590 14720
rect 50270 14655 50590 14656
rect 4190 14176 4510 14177
rect 4190 14112 4198 14176
rect 4262 14112 4278 14176
rect 4342 14112 4358 14176
rect 4422 14112 4438 14176
rect 4502 14112 4510 14176
rect 4190 14111 4510 14112
rect 34910 14176 35230 14177
rect 34910 14112 34918 14176
rect 34982 14112 34998 14176
rect 35062 14112 35078 14176
rect 35142 14112 35158 14176
rect 35222 14112 35230 14176
rect 34910 14111 35230 14112
rect 7999 13834 8065 13837
rect 12507 13834 12573 13837
rect 7999 13832 12573 13834
rect 7999 13776 8004 13832
rect 8060 13776 12512 13832
rect 12568 13776 12573 13832
rect 7999 13774 12573 13776
rect 7999 13771 8065 13774
rect 12507 13771 12573 13774
rect 19550 13632 19870 13633
rect 19550 13568 19558 13632
rect 19622 13568 19638 13632
rect 19702 13568 19718 13632
rect 19782 13568 19798 13632
rect 19862 13568 19870 13632
rect 19550 13567 19870 13568
rect 50270 13632 50590 13633
rect 50270 13568 50278 13632
rect 50342 13568 50358 13632
rect 50422 13568 50438 13632
rect 50502 13568 50518 13632
rect 50582 13568 50590 13632
rect 50270 13567 50590 13568
rect 4190 13088 4510 13089
rect 4190 13024 4198 13088
rect 4262 13024 4278 13088
rect 4342 13024 4358 13088
rect 4422 13024 4438 13088
rect 4502 13024 4510 13088
rect 4190 13023 4510 13024
rect 34910 13088 35230 13089
rect 34910 13024 34918 13088
rect 34982 13024 34998 13088
rect 35062 13024 35078 13088
rect 35142 13024 35158 13088
rect 35222 13024 35230 13088
rect 34910 13023 35230 13024
rect 19550 12544 19870 12545
rect 19550 12480 19558 12544
rect 19622 12480 19638 12544
rect 19702 12480 19718 12544
rect 19782 12480 19798 12544
rect 19862 12480 19870 12544
rect 19550 12479 19870 12480
rect 50270 12544 50590 12545
rect 50270 12480 50278 12544
rect 50342 12480 50358 12544
rect 50422 12480 50438 12544
rect 50502 12480 50518 12544
rect 50582 12480 50590 12544
rect 50270 12479 50590 12480
rect 5791 12066 5857 12069
rect 6803 12066 6869 12069
rect 5791 12064 6869 12066
rect 5791 12008 5796 12064
rect 5852 12008 6808 12064
rect 6864 12008 6869 12064
rect 5791 12006 6869 12008
rect 5791 12003 5857 12006
rect 6803 12003 6869 12006
rect 4190 12000 4510 12001
rect 4190 11936 4198 12000
rect 4262 11936 4278 12000
rect 4342 11936 4358 12000
rect 4422 11936 4438 12000
rect 4502 11936 4510 12000
rect 4190 11935 4510 11936
rect 34910 12000 35230 12001
rect 34910 11936 34918 12000
rect 34982 11936 34998 12000
rect 35062 11936 35078 12000
rect 35142 11936 35158 12000
rect 35222 11936 35230 12000
rect 34910 11935 35230 11936
rect 8091 11794 8157 11797
rect 11679 11794 11745 11797
rect 8091 11792 11745 11794
rect 8091 11736 8096 11792
rect 8152 11736 11684 11792
rect 11740 11736 11745 11792
rect 8091 11734 11745 11736
rect 8091 11731 8157 11734
rect 11679 11731 11745 11734
rect 15175 11794 15241 11797
rect 15175 11792 15376 11794
rect 15175 11736 15180 11792
rect 15236 11736 15376 11792
rect 15175 11734 15376 11736
rect 15175 11731 15241 11734
rect 15316 11658 15376 11734
rect 24743 11658 24809 11661
rect 15316 11656 24809 11658
rect 15316 11600 24748 11656
rect 24804 11600 24809 11656
rect 15316 11598 24809 11600
rect 24743 11595 24809 11598
rect 19550 11456 19870 11457
rect 19550 11392 19558 11456
rect 19622 11392 19638 11456
rect 19702 11392 19718 11456
rect 19782 11392 19798 11456
rect 19862 11392 19870 11456
rect 19550 11391 19870 11392
rect 50270 11456 50590 11457
rect 50270 11392 50278 11456
rect 50342 11392 50358 11456
rect 50422 11392 50438 11456
rect 50502 11392 50518 11456
rect 50582 11392 50590 11456
rect 50270 11391 50590 11392
rect 4190 10912 4510 10913
rect 4190 10848 4198 10912
rect 4262 10848 4278 10912
rect 4342 10848 4358 10912
rect 4422 10848 4438 10912
rect 4502 10848 4510 10912
rect 4190 10847 4510 10848
rect 34910 10912 35230 10913
rect 34910 10848 34918 10912
rect 34982 10848 34998 10912
rect 35062 10848 35078 10912
rect 35142 10848 35158 10912
rect 35222 10848 35230 10912
rect 34910 10847 35230 10848
rect 19550 10368 19870 10369
rect 19550 10304 19558 10368
rect 19622 10304 19638 10368
rect 19702 10304 19718 10368
rect 19782 10304 19798 10368
rect 19862 10304 19870 10368
rect 19550 10303 19870 10304
rect 50270 10368 50590 10369
rect 50270 10304 50278 10368
rect 50342 10304 50358 10368
rect 50422 10304 50438 10368
rect 50502 10304 50518 10368
rect 50582 10304 50590 10368
rect 50270 10303 50590 10304
rect 4190 9824 4510 9825
rect 4190 9760 4198 9824
rect 4262 9760 4278 9824
rect 4342 9760 4358 9824
rect 4422 9760 4438 9824
rect 4502 9760 4510 9824
rect 4190 9759 4510 9760
rect 34910 9824 35230 9825
rect 34910 9760 34918 9824
rect 34982 9760 34998 9824
rect 35062 9760 35078 9824
rect 35142 9760 35158 9824
rect 35222 9760 35230 9824
rect 34910 9759 35230 9760
rect 49215 9618 49281 9621
rect 57127 9618 57193 9621
rect 49215 9616 57193 9618
rect 49215 9560 49220 9616
rect 49276 9560 57132 9616
rect 57188 9560 57193 9616
rect 49215 9558 57193 9560
rect 49215 9555 49281 9558
rect 57127 9555 57193 9558
rect 19550 9280 19870 9281
rect 19550 9216 19558 9280
rect 19622 9216 19638 9280
rect 19702 9216 19718 9280
rect 19782 9216 19798 9280
rect 19862 9216 19870 9280
rect 19550 9215 19870 9216
rect 50270 9280 50590 9281
rect 50270 9216 50278 9280
rect 50342 9216 50358 9280
rect 50422 9216 50438 9280
rect 50502 9216 50518 9280
rect 50582 9216 50590 9280
rect 50270 9215 50590 9216
rect 4190 8736 4510 8737
rect 4190 8672 4198 8736
rect 4262 8672 4278 8736
rect 4342 8672 4358 8736
rect 4422 8672 4438 8736
rect 4502 8672 4510 8736
rect 4190 8671 4510 8672
rect 34910 8736 35230 8737
rect 34910 8672 34918 8736
rect 34982 8672 34998 8736
rect 35062 8672 35078 8736
rect 35142 8672 35158 8736
rect 35222 8672 35230 8736
rect 34910 8671 35230 8672
rect 19550 8192 19870 8193
rect 19550 8128 19558 8192
rect 19622 8128 19638 8192
rect 19702 8128 19718 8192
rect 19782 8128 19798 8192
rect 19862 8128 19870 8192
rect 19550 8127 19870 8128
rect 50270 8192 50590 8193
rect 50270 8128 50278 8192
rect 50342 8128 50358 8192
rect 50422 8128 50438 8192
rect 50502 8128 50518 8192
rect 50582 8128 50590 8192
rect 50270 8127 50590 8128
rect 19867 7714 19933 7717
rect 20276 7714 20282 7716
rect 19867 7712 20282 7714
rect 19867 7656 19872 7712
rect 19928 7656 20282 7712
rect 19867 7654 20282 7656
rect 19867 7651 19933 7654
rect 20276 7652 20282 7654
rect 20346 7652 20352 7716
rect 4190 7648 4510 7649
rect 4190 7584 4198 7648
rect 4262 7584 4278 7648
rect 4342 7584 4358 7648
rect 4422 7584 4438 7648
rect 4502 7584 4510 7648
rect 4190 7583 4510 7584
rect 34910 7648 35230 7649
rect 34910 7584 34918 7648
rect 34982 7584 34998 7648
rect 35062 7584 35078 7648
rect 35142 7584 35158 7648
rect 35222 7584 35230 7648
rect 34910 7583 35230 7584
rect 19867 7578 19933 7581
rect 20143 7578 20209 7581
rect 19867 7576 20209 7578
rect 19867 7520 19872 7576
rect 19928 7520 20148 7576
rect 20204 7520 20209 7576
rect 19867 7518 20209 7520
rect 19867 7515 19933 7518
rect 20143 7515 20209 7518
rect 19550 7104 19870 7105
rect 19550 7040 19558 7104
rect 19622 7040 19638 7104
rect 19702 7040 19718 7104
rect 19782 7040 19798 7104
rect 19862 7040 19870 7104
rect 19550 7039 19870 7040
rect 50270 7104 50590 7105
rect 50270 7040 50278 7104
rect 50342 7040 50358 7104
rect 50422 7040 50438 7104
rect 50502 7040 50518 7104
rect 50582 7040 50590 7104
rect 50270 7039 50590 7040
rect 4190 6560 4510 6561
rect 4190 6496 4198 6560
rect 4262 6496 4278 6560
rect 4342 6496 4358 6560
rect 4422 6496 4438 6560
rect 4502 6496 4510 6560
rect 4190 6495 4510 6496
rect 34910 6560 35230 6561
rect 34910 6496 34918 6560
rect 34982 6496 34998 6560
rect 35062 6496 35078 6560
rect 35142 6496 35158 6560
rect 35222 6496 35230 6560
rect 34910 6495 35230 6496
rect 19550 6016 19870 6017
rect 19550 5952 19558 6016
rect 19622 5952 19638 6016
rect 19702 5952 19718 6016
rect 19782 5952 19798 6016
rect 19862 5952 19870 6016
rect 19550 5951 19870 5952
rect 50270 6016 50590 6017
rect 50270 5952 50278 6016
rect 50342 5952 50358 6016
rect 50422 5952 50438 6016
rect 50502 5952 50518 6016
rect 50582 5952 50590 6016
rect 50270 5951 50590 5952
rect 4190 5472 4510 5473
rect 4190 5408 4198 5472
rect 4262 5408 4278 5472
rect 4342 5408 4358 5472
rect 4422 5408 4438 5472
rect 4502 5408 4510 5472
rect 4190 5407 4510 5408
rect 34910 5472 35230 5473
rect 34910 5408 34918 5472
rect 34982 5408 34998 5472
rect 35062 5408 35078 5472
rect 35142 5408 35158 5472
rect 35222 5408 35230 5472
rect 34910 5407 35230 5408
rect 19550 4928 19870 4929
rect 19550 4864 19558 4928
rect 19622 4864 19638 4928
rect 19702 4864 19718 4928
rect 19782 4864 19798 4928
rect 19862 4864 19870 4928
rect 19550 4863 19870 4864
rect 50270 4928 50590 4929
rect 50270 4864 50278 4928
rect 50342 4864 50358 4928
rect 50422 4864 50438 4928
rect 50502 4864 50518 4928
rect 50582 4864 50590 4928
rect 50270 4863 50590 4864
rect 4190 4384 4510 4385
rect 4190 4320 4198 4384
rect 4262 4320 4278 4384
rect 4342 4320 4358 4384
rect 4422 4320 4438 4384
rect 4502 4320 4510 4384
rect 4190 4319 4510 4320
rect 34910 4384 35230 4385
rect 34910 4320 34918 4384
rect 34982 4320 34998 4384
rect 35062 4320 35078 4384
rect 35142 4320 35158 4384
rect 35222 4320 35230 4384
rect 34910 4319 35230 4320
rect 7723 4042 7789 4045
rect 43511 4042 43577 4045
rect 7723 4040 43577 4042
rect 7723 3984 7728 4040
rect 7784 3984 43516 4040
rect 43572 3984 43577 4040
rect 7723 3982 43577 3984
rect 7723 3979 7789 3982
rect 43511 3979 43577 3982
rect 31735 3906 31801 3909
rect 33023 3906 33089 3909
rect 41252 3906 41258 3908
rect 31735 3904 33089 3906
rect 31735 3848 31740 3904
rect 31796 3848 33028 3904
rect 33084 3848 33089 3904
rect 31735 3846 33089 3848
rect 31735 3843 31801 3846
rect 33023 3843 33089 3846
rect 33164 3846 41258 3906
rect 19550 3840 19870 3841
rect 19550 3776 19558 3840
rect 19622 3776 19638 3840
rect 19702 3776 19718 3840
rect 19782 3776 19798 3840
rect 19862 3776 19870 3840
rect 19550 3775 19870 3776
rect 14347 3770 14413 3773
rect 18947 3770 19013 3773
rect 14347 3768 19013 3770
rect 14347 3712 14352 3768
rect 14408 3712 18952 3768
rect 19008 3712 19013 3768
rect 14347 3710 19013 3712
rect 14347 3707 14413 3710
rect 18947 3707 19013 3710
rect 32471 3770 32537 3773
rect 33164 3770 33224 3846
rect 41252 3844 41258 3846
rect 41322 3844 41328 3908
rect 50270 3840 50590 3841
rect 50270 3776 50278 3840
rect 50342 3776 50358 3840
rect 50422 3776 50438 3840
rect 50502 3776 50518 3840
rect 50582 3776 50590 3840
rect 50270 3775 50590 3776
rect 32471 3768 33224 3770
rect 32471 3712 32476 3768
rect 32532 3712 33224 3768
rect 32471 3710 33224 3712
rect 34035 3770 34101 3773
rect 44615 3770 44681 3773
rect 34035 3768 44681 3770
rect 34035 3712 34040 3768
rect 34096 3712 44620 3768
rect 44676 3712 44681 3768
rect 34035 3710 44681 3712
rect 32471 3707 32537 3710
rect 34035 3707 34101 3710
rect 44615 3707 44681 3710
rect 11127 3634 11193 3637
rect 47191 3634 47257 3637
rect 11127 3632 47257 3634
rect 11127 3576 11132 3632
rect 11188 3576 47196 3632
rect 47252 3576 47257 3632
rect 11127 3574 47257 3576
rect 11127 3571 11193 3574
rect 47191 3571 47257 3574
rect 11219 3498 11285 3501
rect 11219 3496 48496 3498
rect 11219 3440 11224 3496
rect 11280 3440 48496 3496
rect 11219 3438 48496 3440
rect 11219 3435 11285 3438
rect 48436 3365 48496 3438
rect 18119 3362 18185 3365
rect 26859 3362 26925 3365
rect 18119 3360 26925 3362
rect 18119 3304 18124 3360
rect 18180 3304 26864 3360
rect 26920 3304 26925 3360
rect 18119 3302 26925 3304
rect 18119 3299 18185 3302
rect 26859 3299 26925 3302
rect 31827 3362 31893 3365
rect 33667 3362 33733 3365
rect 31827 3360 33733 3362
rect 31827 3304 31832 3360
rect 31888 3304 33672 3360
rect 33728 3304 33733 3360
rect 31827 3302 33733 3304
rect 31827 3299 31893 3302
rect 33667 3299 33733 3302
rect 48387 3360 48496 3365
rect 48387 3304 48392 3360
rect 48448 3304 48496 3360
rect 48387 3302 48496 3304
rect 48387 3299 48453 3302
rect 4190 3296 4510 3297
rect 4190 3232 4198 3296
rect 4262 3232 4278 3296
rect 4342 3232 4358 3296
rect 4422 3232 4438 3296
rect 4502 3232 4510 3296
rect 4190 3231 4510 3232
rect 34910 3296 35230 3297
rect 34910 3232 34918 3296
rect 34982 3232 34998 3296
rect 35062 3232 35078 3296
rect 35142 3232 35158 3296
rect 35222 3232 35230 3296
rect 34910 3231 35230 3232
rect 18211 3226 18277 3229
rect 34495 3226 34561 3229
rect 18211 3224 34561 3226
rect 18211 3168 18216 3224
rect 18272 3168 34500 3224
rect 34556 3168 34561 3224
rect 18211 3166 34561 3168
rect 18211 3163 18277 3166
rect 34495 3163 34561 3166
rect 9195 3090 9261 3093
rect 42039 3090 42105 3093
rect 9195 3088 42105 3090
rect 9195 3032 9200 3088
rect 9256 3032 42044 3088
rect 42100 3032 42105 3088
rect 9195 3030 42105 3032
rect 9195 3027 9261 3030
rect 42039 3027 42105 3030
rect 34495 2954 34561 2957
rect 35415 2954 35481 2957
rect 34495 2952 35481 2954
rect 34495 2896 34500 2952
rect 34556 2896 35420 2952
rect 35476 2896 35481 2952
rect 34495 2894 35481 2896
rect 34495 2891 34561 2894
rect 35415 2891 35481 2894
rect 38635 2954 38701 2957
rect 41119 2954 41185 2957
rect 38635 2952 41185 2954
rect 38635 2896 38640 2952
rect 38696 2896 41124 2952
rect 41180 2896 41185 2952
rect 38635 2894 41185 2896
rect 38635 2891 38701 2894
rect 41119 2891 41185 2894
rect 41252 2892 41258 2956
rect 41322 2954 41328 2956
rect 55655 2954 55721 2957
rect 41322 2952 55721 2954
rect 41322 2896 55660 2952
rect 55716 2896 55721 2952
rect 41322 2894 55721 2896
rect 41322 2892 41328 2894
rect 55655 2891 55721 2894
rect 26859 2818 26925 2821
rect 37623 2818 37689 2821
rect 26859 2816 37689 2818
rect 26859 2760 26864 2816
rect 26920 2760 37628 2816
rect 37684 2760 37689 2816
rect 26859 2758 37689 2760
rect 26859 2755 26925 2758
rect 37623 2755 37689 2758
rect 19550 2752 19870 2753
rect 19550 2688 19558 2752
rect 19622 2688 19638 2752
rect 19702 2688 19718 2752
rect 19782 2688 19798 2752
rect 19862 2688 19870 2752
rect 19550 2687 19870 2688
rect 50270 2752 50590 2753
rect 50270 2688 50278 2752
rect 50342 2688 50358 2752
rect 50422 2688 50438 2752
rect 50502 2688 50518 2752
rect 50582 2688 50590 2752
rect 50270 2687 50590 2688
rect 4190 2208 4510 2209
rect 4190 2144 4198 2208
rect 4262 2144 4278 2208
rect 4342 2144 4358 2208
rect 4422 2144 4438 2208
rect 4502 2144 4510 2208
rect 4190 2143 4510 2144
rect 34910 2208 35230 2209
rect 34910 2144 34918 2208
rect 34982 2144 34998 2208
rect 35062 2144 35078 2208
rect 35142 2144 35158 2208
rect 35222 2144 35230 2208
rect 34910 2143 35230 2144
rect 20276 852 20282 916
rect 20346 914 20352 916
rect 20419 914 20485 917
rect 20346 912 20485 914
rect 20346 856 20424 912
rect 20480 856 20485 912
rect 20346 854 20485 856
rect 20346 852 20352 854
rect 20419 851 20485 854
<< via3 >>
rect 4198 57692 4262 57696
rect 4198 57636 4202 57692
rect 4202 57636 4258 57692
rect 4258 57636 4262 57692
rect 4198 57632 4262 57636
rect 4278 57692 4342 57696
rect 4278 57636 4282 57692
rect 4282 57636 4338 57692
rect 4338 57636 4342 57692
rect 4278 57632 4342 57636
rect 4358 57692 4422 57696
rect 4358 57636 4362 57692
rect 4362 57636 4418 57692
rect 4418 57636 4422 57692
rect 4358 57632 4422 57636
rect 4438 57692 4502 57696
rect 4438 57636 4442 57692
rect 4442 57636 4498 57692
rect 4498 57636 4502 57692
rect 4438 57632 4502 57636
rect 34918 57692 34982 57696
rect 34918 57636 34922 57692
rect 34922 57636 34978 57692
rect 34978 57636 34982 57692
rect 34918 57632 34982 57636
rect 34998 57692 35062 57696
rect 34998 57636 35002 57692
rect 35002 57636 35058 57692
rect 35058 57636 35062 57692
rect 34998 57632 35062 57636
rect 35078 57692 35142 57696
rect 35078 57636 35082 57692
rect 35082 57636 35138 57692
rect 35138 57636 35142 57692
rect 35078 57632 35142 57636
rect 35158 57692 35222 57696
rect 35158 57636 35162 57692
rect 35162 57636 35218 57692
rect 35218 57636 35222 57692
rect 35158 57632 35222 57636
rect 19558 57148 19622 57152
rect 19558 57092 19562 57148
rect 19562 57092 19618 57148
rect 19618 57092 19622 57148
rect 19558 57088 19622 57092
rect 19638 57148 19702 57152
rect 19638 57092 19642 57148
rect 19642 57092 19698 57148
rect 19698 57092 19702 57148
rect 19638 57088 19702 57092
rect 19718 57148 19782 57152
rect 19718 57092 19722 57148
rect 19722 57092 19778 57148
rect 19778 57092 19782 57148
rect 19718 57088 19782 57092
rect 19798 57148 19862 57152
rect 19798 57092 19802 57148
rect 19802 57092 19858 57148
rect 19858 57092 19862 57148
rect 19798 57088 19862 57092
rect 50278 57148 50342 57152
rect 50278 57092 50282 57148
rect 50282 57092 50338 57148
rect 50338 57092 50342 57148
rect 50278 57088 50342 57092
rect 50358 57148 50422 57152
rect 50358 57092 50362 57148
rect 50362 57092 50418 57148
rect 50418 57092 50422 57148
rect 50358 57088 50422 57092
rect 50438 57148 50502 57152
rect 50438 57092 50442 57148
rect 50442 57092 50498 57148
rect 50498 57092 50502 57148
rect 50438 57088 50502 57092
rect 50518 57148 50582 57152
rect 50518 57092 50522 57148
rect 50522 57092 50578 57148
rect 50578 57092 50582 57148
rect 50518 57088 50582 57092
rect 4198 56604 4262 56608
rect 4198 56548 4202 56604
rect 4202 56548 4258 56604
rect 4258 56548 4262 56604
rect 4198 56544 4262 56548
rect 4278 56604 4342 56608
rect 4278 56548 4282 56604
rect 4282 56548 4338 56604
rect 4338 56548 4342 56604
rect 4278 56544 4342 56548
rect 4358 56604 4422 56608
rect 4358 56548 4362 56604
rect 4362 56548 4418 56604
rect 4418 56548 4422 56604
rect 4358 56544 4422 56548
rect 4438 56604 4502 56608
rect 4438 56548 4442 56604
rect 4442 56548 4498 56604
rect 4498 56548 4502 56604
rect 4438 56544 4502 56548
rect 34918 56604 34982 56608
rect 34918 56548 34922 56604
rect 34922 56548 34978 56604
rect 34978 56548 34982 56604
rect 34918 56544 34982 56548
rect 34998 56604 35062 56608
rect 34998 56548 35002 56604
rect 35002 56548 35058 56604
rect 35058 56548 35062 56604
rect 34998 56544 35062 56548
rect 35078 56604 35142 56608
rect 35078 56548 35082 56604
rect 35082 56548 35138 56604
rect 35138 56548 35142 56604
rect 35078 56544 35142 56548
rect 35158 56604 35222 56608
rect 35158 56548 35162 56604
rect 35162 56548 35218 56604
rect 35218 56548 35222 56604
rect 35158 56544 35222 56548
rect 19558 56060 19622 56064
rect 19558 56004 19562 56060
rect 19562 56004 19618 56060
rect 19618 56004 19622 56060
rect 19558 56000 19622 56004
rect 19638 56060 19702 56064
rect 19638 56004 19642 56060
rect 19642 56004 19698 56060
rect 19698 56004 19702 56060
rect 19638 56000 19702 56004
rect 19718 56060 19782 56064
rect 19718 56004 19722 56060
rect 19722 56004 19778 56060
rect 19778 56004 19782 56060
rect 19718 56000 19782 56004
rect 19798 56060 19862 56064
rect 19798 56004 19802 56060
rect 19802 56004 19858 56060
rect 19858 56004 19862 56060
rect 19798 56000 19862 56004
rect 50278 56060 50342 56064
rect 50278 56004 50282 56060
rect 50282 56004 50338 56060
rect 50338 56004 50342 56060
rect 50278 56000 50342 56004
rect 50358 56060 50422 56064
rect 50358 56004 50362 56060
rect 50362 56004 50418 56060
rect 50418 56004 50422 56060
rect 50358 56000 50422 56004
rect 50438 56060 50502 56064
rect 50438 56004 50442 56060
rect 50442 56004 50498 56060
rect 50498 56004 50502 56060
rect 50438 56000 50502 56004
rect 50518 56060 50582 56064
rect 50518 56004 50522 56060
rect 50522 56004 50578 56060
rect 50578 56004 50582 56060
rect 50518 56000 50582 56004
rect 4198 55516 4262 55520
rect 4198 55460 4202 55516
rect 4202 55460 4258 55516
rect 4258 55460 4262 55516
rect 4198 55456 4262 55460
rect 4278 55516 4342 55520
rect 4278 55460 4282 55516
rect 4282 55460 4338 55516
rect 4338 55460 4342 55516
rect 4278 55456 4342 55460
rect 4358 55516 4422 55520
rect 4358 55460 4362 55516
rect 4362 55460 4418 55516
rect 4418 55460 4422 55516
rect 4358 55456 4422 55460
rect 4438 55516 4502 55520
rect 4438 55460 4442 55516
rect 4442 55460 4498 55516
rect 4498 55460 4502 55516
rect 4438 55456 4502 55460
rect 34918 55516 34982 55520
rect 34918 55460 34922 55516
rect 34922 55460 34978 55516
rect 34978 55460 34982 55516
rect 34918 55456 34982 55460
rect 34998 55516 35062 55520
rect 34998 55460 35002 55516
rect 35002 55460 35058 55516
rect 35058 55460 35062 55516
rect 34998 55456 35062 55460
rect 35078 55516 35142 55520
rect 35078 55460 35082 55516
rect 35082 55460 35138 55516
rect 35138 55460 35142 55516
rect 35078 55456 35142 55460
rect 35158 55516 35222 55520
rect 35158 55460 35162 55516
rect 35162 55460 35218 55516
rect 35218 55460 35222 55516
rect 35158 55456 35222 55460
rect 19558 54972 19622 54976
rect 19558 54916 19562 54972
rect 19562 54916 19618 54972
rect 19618 54916 19622 54972
rect 19558 54912 19622 54916
rect 19638 54972 19702 54976
rect 19638 54916 19642 54972
rect 19642 54916 19698 54972
rect 19698 54916 19702 54972
rect 19638 54912 19702 54916
rect 19718 54972 19782 54976
rect 19718 54916 19722 54972
rect 19722 54916 19778 54972
rect 19778 54916 19782 54972
rect 19718 54912 19782 54916
rect 19798 54972 19862 54976
rect 19798 54916 19802 54972
rect 19802 54916 19858 54972
rect 19858 54916 19862 54972
rect 19798 54912 19862 54916
rect 50278 54972 50342 54976
rect 50278 54916 50282 54972
rect 50282 54916 50338 54972
rect 50338 54916 50342 54972
rect 50278 54912 50342 54916
rect 50358 54972 50422 54976
rect 50358 54916 50362 54972
rect 50362 54916 50418 54972
rect 50418 54916 50422 54972
rect 50358 54912 50422 54916
rect 50438 54972 50502 54976
rect 50438 54916 50442 54972
rect 50442 54916 50498 54972
rect 50498 54916 50502 54972
rect 50438 54912 50502 54916
rect 50518 54972 50582 54976
rect 50518 54916 50522 54972
rect 50522 54916 50578 54972
rect 50578 54916 50582 54972
rect 50518 54912 50582 54916
rect 4198 54428 4262 54432
rect 4198 54372 4202 54428
rect 4202 54372 4258 54428
rect 4258 54372 4262 54428
rect 4198 54368 4262 54372
rect 4278 54428 4342 54432
rect 4278 54372 4282 54428
rect 4282 54372 4338 54428
rect 4338 54372 4342 54428
rect 4278 54368 4342 54372
rect 4358 54428 4422 54432
rect 4358 54372 4362 54428
rect 4362 54372 4418 54428
rect 4418 54372 4422 54428
rect 4358 54368 4422 54372
rect 4438 54428 4502 54432
rect 4438 54372 4442 54428
rect 4442 54372 4498 54428
rect 4498 54372 4502 54428
rect 4438 54368 4502 54372
rect 34918 54428 34982 54432
rect 34918 54372 34922 54428
rect 34922 54372 34978 54428
rect 34978 54372 34982 54428
rect 34918 54368 34982 54372
rect 34998 54428 35062 54432
rect 34998 54372 35002 54428
rect 35002 54372 35058 54428
rect 35058 54372 35062 54428
rect 34998 54368 35062 54372
rect 35078 54428 35142 54432
rect 35078 54372 35082 54428
rect 35082 54372 35138 54428
rect 35138 54372 35142 54428
rect 35078 54368 35142 54372
rect 35158 54428 35222 54432
rect 35158 54372 35162 54428
rect 35162 54372 35218 54428
rect 35218 54372 35222 54428
rect 35158 54368 35222 54372
rect 19558 53884 19622 53888
rect 19558 53828 19562 53884
rect 19562 53828 19618 53884
rect 19618 53828 19622 53884
rect 19558 53824 19622 53828
rect 19638 53884 19702 53888
rect 19638 53828 19642 53884
rect 19642 53828 19698 53884
rect 19698 53828 19702 53884
rect 19638 53824 19702 53828
rect 19718 53884 19782 53888
rect 19718 53828 19722 53884
rect 19722 53828 19778 53884
rect 19778 53828 19782 53884
rect 19718 53824 19782 53828
rect 19798 53884 19862 53888
rect 19798 53828 19802 53884
rect 19802 53828 19858 53884
rect 19858 53828 19862 53884
rect 19798 53824 19862 53828
rect 50278 53884 50342 53888
rect 50278 53828 50282 53884
rect 50282 53828 50338 53884
rect 50338 53828 50342 53884
rect 50278 53824 50342 53828
rect 50358 53884 50422 53888
rect 50358 53828 50362 53884
rect 50362 53828 50418 53884
rect 50418 53828 50422 53884
rect 50358 53824 50422 53828
rect 50438 53884 50502 53888
rect 50438 53828 50442 53884
rect 50442 53828 50498 53884
rect 50498 53828 50502 53884
rect 50438 53824 50502 53828
rect 50518 53884 50582 53888
rect 50518 53828 50522 53884
rect 50522 53828 50578 53884
rect 50578 53828 50582 53884
rect 50518 53824 50582 53828
rect 4198 53340 4262 53344
rect 4198 53284 4202 53340
rect 4202 53284 4258 53340
rect 4258 53284 4262 53340
rect 4198 53280 4262 53284
rect 4278 53340 4342 53344
rect 4278 53284 4282 53340
rect 4282 53284 4338 53340
rect 4338 53284 4342 53340
rect 4278 53280 4342 53284
rect 4358 53340 4422 53344
rect 4358 53284 4362 53340
rect 4362 53284 4418 53340
rect 4418 53284 4422 53340
rect 4358 53280 4422 53284
rect 4438 53340 4502 53344
rect 4438 53284 4442 53340
rect 4442 53284 4498 53340
rect 4498 53284 4502 53340
rect 4438 53280 4502 53284
rect 34918 53340 34982 53344
rect 34918 53284 34922 53340
rect 34922 53284 34978 53340
rect 34978 53284 34982 53340
rect 34918 53280 34982 53284
rect 34998 53340 35062 53344
rect 34998 53284 35002 53340
rect 35002 53284 35058 53340
rect 35058 53284 35062 53340
rect 34998 53280 35062 53284
rect 35078 53340 35142 53344
rect 35078 53284 35082 53340
rect 35082 53284 35138 53340
rect 35138 53284 35142 53340
rect 35078 53280 35142 53284
rect 35158 53340 35222 53344
rect 35158 53284 35162 53340
rect 35162 53284 35218 53340
rect 35218 53284 35222 53340
rect 35158 53280 35222 53284
rect 19558 52796 19622 52800
rect 19558 52740 19562 52796
rect 19562 52740 19618 52796
rect 19618 52740 19622 52796
rect 19558 52736 19622 52740
rect 19638 52796 19702 52800
rect 19638 52740 19642 52796
rect 19642 52740 19698 52796
rect 19698 52740 19702 52796
rect 19638 52736 19702 52740
rect 19718 52796 19782 52800
rect 19718 52740 19722 52796
rect 19722 52740 19778 52796
rect 19778 52740 19782 52796
rect 19718 52736 19782 52740
rect 19798 52796 19862 52800
rect 19798 52740 19802 52796
rect 19802 52740 19858 52796
rect 19858 52740 19862 52796
rect 19798 52736 19862 52740
rect 50278 52796 50342 52800
rect 50278 52740 50282 52796
rect 50282 52740 50338 52796
rect 50338 52740 50342 52796
rect 50278 52736 50342 52740
rect 50358 52796 50422 52800
rect 50358 52740 50362 52796
rect 50362 52740 50418 52796
rect 50418 52740 50422 52796
rect 50358 52736 50422 52740
rect 50438 52796 50502 52800
rect 50438 52740 50442 52796
rect 50442 52740 50498 52796
rect 50498 52740 50502 52796
rect 50438 52736 50502 52740
rect 50518 52796 50582 52800
rect 50518 52740 50522 52796
rect 50522 52740 50578 52796
rect 50578 52740 50582 52796
rect 50518 52736 50582 52740
rect 4198 52252 4262 52256
rect 4198 52196 4202 52252
rect 4202 52196 4258 52252
rect 4258 52196 4262 52252
rect 4198 52192 4262 52196
rect 4278 52252 4342 52256
rect 4278 52196 4282 52252
rect 4282 52196 4338 52252
rect 4338 52196 4342 52252
rect 4278 52192 4342 52196
rect 4358 52252 4422 52256
rect 4358 52196 4362 52252
rect 4362 52196 4418 52252
rect 4418 52196 4422 52252
rect 4358 52192 4422 52196
rect 4438 52252 4502 52256
rect 4438 52196 4442 52252
rect 4442 52196 4498 52252
rect 4498 52196 4502 52252
rect 4438 52192 4502 52196
rect 34918 52252 34982 52256
rect 34918 52196 34922 52252
rect 34922 52196 34978 52252
rect 34978 52196 34982 52252
rect 34918 52192 34982 52196
rect 34998 52252 35062 52256
rect 34998 52196 35002 52252
rect 35002 52196 35058 52252
rect 35058 52196 35062 52252
rect 34998 52192 35062 52196
rect 35078 52252 35142 52256
rect 35078 52196 35082 52252
rect 35082 52196 35138 52252
rect 35138 52196 35142 52252
rect 35078 52192 35142 52196
rect 35158 52252 35222 52256
rect 35158 52196 35162 52252
rect 35162 52196 35218 52252
rect 35218 52196 35222 52252
rect 35158 52192 35222 52196
rect 19558 51708 19622 51712
rect 19558 51652 19562 51708
rect 19562 51652 19618 51708
rect 19618 51652 19622 51708
rect 19558 51648 19622 51652
rect 19638 51708 19702 51712
rect 19638 51652 19642 51708
rect 19642 51652 19698 51708
rect 19698 51652 19702 51708
rect 19638 51648 19702 51652
rect 19718 51708 19782 51712
rect 19718 51652 19722 51708
rect 19722 51652 19778 51708
rect 19778 51652 19782 51708
rect 19718 51648 19782 51652
rect 19798 51708 19862 51712
rect 19798 51652 19802 51708
rect 19802 51652 19858 51708
rect 19858 51652 19862 51708
rect 19798 51648 19862 51652
rect 50278 51708 50342 51712
rect 50278 51652 50282 51708
rect 50282 51652 50338 51708
rect 50338 51652 50342 51708
rect 50278 51648 50342 51652
rect 50358 51708 50422 51712
rect 50358 51652 50362 51708
rect 50362 51652 50418 51708
rect 50418 51652 50422 51708
rect 50358 51648 50422 51652
rect 50438 51708 50502 51712
rect 50438 51652 50442 51708
rect 50442 51652 50498 51708
rect 50498 51652 50502 51708
rect 50438 51648 50502 51652
rect 50518 51708 50582 51712
rect 50518 51652 50522 51708
rect 50522 51652 50578 51708
rect 50578 51652 50582 51708
rect 50518 51648 50582 51652
rect 4198 51164 4262 51168
rect 4198 51108 4202 51164
rect 4202 51108 4258 51164
rect 4258 51108 4262 51164
rect 4198 51104 4262 51108
rect 4278 51164 4342 51168
rect 4278 51108 4282 51164
rect 4282 51108 4338 51164
rect 4338 51108 4342 51164
rect 4278 51104 4342 51108
rect 4358 51164 4422 51168
rect 4358 51108 4362 51164
rect 4362 51108 4418 51164
rect 4418 51108 4422 51164
rect 4358 51104 4422 51108
rect 4438 51164 4502 51168
rect 4438 51108 4442 51164
rect 4442 51108 4498 51164
rect 4498 51108 4502 51164
rect 4438 51104 4502 51108
rect 34918 51164 34982 51168
rect 34918 51108 34922 51164
rect 34922 51108 34978 51164
rect 34978 51108 34982 51164
rect 34918 51104 34982 51108
rect 34998 51164 35062 51168
rect 34998 51108 35002 51164
rect 35002 51108 35058 51164
rect 35058 51108 35062 51164
rect 34998 51104 35062 51108
rect 35078 51164 35142 51168
rect 35078 51108 35082 51164
rect 35082 51108 35138 51164
rect 35138 51108 35142 51164
rect 35078 51104 35142 51108
rect 35158 51164 35222 51168
rect 35158 51108 35162 51164
rect 35162 51108 35218 51164
rect 35218 51108 35222 51164
rect 35158 51104 35222 51108
rect 19558 50620 19622 50624
rect 19558 50564 19562 50620
rect 19562 50564 19618 50620
rect 19618 50564 19622 50620
rect 19558 50560 19622 50564
rect 19638 50620 19702 50624
rect 19638 50564 19642 50620
rect 19642 50564 19698 50620
rect 19698 50564 19702 50620
rect 19638 50560 19702 50564
rect 19718 50620 19782 50624
rect 19718 50564 19722 50620
rect 19722 50564 19778 50620
rect 19778 50564 19782 50620
rect 19718 50560 19782 50564
rect 19798 50620 19862 50624
rect 19798 50564 19802 50620
rect 19802 50564 19858 50620
rect 19858 50564 19862 50620
rect 19798 50560 19862 50564
rect 50278 50620 50342 50624
rect 50278 50564 50282 50620
rect 50282 50564 50338 50620
rect 50338 50564 50342 50620
rect 50278 50560 50342 50564
rect 50358 50620 50422 50624
rect 50358 50564 50362 50620
rect 50362 50564 50418 50620
rect 50418 50564 50422 50620
rect 50358 50560 50422 50564
rect 50438 50620 50502 50624
rect 50438 50564 50442 50620
rect 50442 50564 50498 50620
rect 50498 50564 50502 50620
rect 50438 50560 50502 50564
rect 50518 50620 50582 50624
rect 50518 50564 50522 50620
rect 50522 50564 50578 50620
rect 50578 50564 50582 50620
rect 50518 50560 50582 50564
rect 4198 50076 4262 50080
rect 4198 50020 4202 50076
rect 4202 50020 4258 50076
rect 4258 50020 4262 50076
rect 4198 50016 4262 50020
rect 4278 50076 4342 50080
rect 4278 50020 4282 50076
rect 4282 50020 4338 50076
rect 4338 50020 4342 50076
rect 4278 50016 4342 50020
rect 4358 50076 4422 50080
rect 4358 50020 4362 50076
rect 4362 50020 4418 50076
rect 4418 50020 4422 50076
rect 4358 50016 4422 50020
rect 4438 50076 4502 50080
rect 4438 50020 4442 50076
rect 4442 50020 4498 50076
rect 4498 50020 4502 50076
rect 4438 50016 4502 50020
rect 34918 50076 34982 50080
rect 34918 50020 34922 50076
rect 34922 50020 34978 50076
rect 34978 50020 34982 50076
rect 34918 50016 34982 50020
rect 34998 50076 35062 50080
rect 34998 50020 35002 50076
rect 35002 50020 35058 50076
rect 35058 50020 35062 50076
rect 34998 50016 35062 50020
rect 35078 50076 35142 50080
rect 35078 50020 35082 50076
rect 35082 50020 35138 50076
rect 35138 50020 35142 50076
rect 35078 50016 35142 50020
rect 35158 50076 35222 50080
rect 35158 50020 35162 50076
rect 35162 50020 35218 50076
rect 35218 50020 35222 50076
rect 35158 50016 35222 50020
rect 19558 49532 19622 49536
rect 19558 49476 19562 49532
rect 19562 49476 19618 49532
rect 19618 49476 19622 49532
rect 19558 49472 19622 49476
rect 19638 49532 19702 49536
rect 19638 49476 19642 49532
rect 19642 49476 19698 49532
rect 19698 49476 19702 49532
rect 19638 49472 19702 49476
rect 19718 49532 19782 49536
rect 19718 49476 19722 49532
rect 19722 49476 19778 49532
rect 19778 49476 19782 49532
rect 19718 49472 19782 49476
rect 19798 49532 19862 49536
rect 19798 49476 19802 49532
rect 19802 49476 19858 49532
rect 19858 49476 19862 49532
rect 19798 49472 19862 49476
rect 50278 49532 50342 49536
rect 50278 49476 50282 49532
rect 50282 49476 50338 49532
rect 50338 49476 50342 49532
rect 50278 49472 50342 49476
rect 50358 49532 50422 49536
rect 50358 49476 50362 49532
rect 50362 49476 50418 49532
rect 50418 49476 50422 49532
rect 50358 49472 50422 49476
rect 50438 49532 50502 49536
rect 50438 49476 50442 49532
rect 50442 49476 50498 49532
rect 50498 49476 50502 49532
rect 50438 49472 50502 49476
rect 50518 49532 50582 49536
rect 50518 49476 50522 49532
rect 50522 49476 50578 49532
rect 50578 49476 50582 49532
rect 50518 49472 50582 49476
rect 4198 48988 4262 48992
rect 4198 48932 4202 48988
rect 4202 48932 4258 48988
rect 4258 48932 4262 48988
rect 4198 48928 4262 48932
rect 4278 48988 4342 48992
rect 4278 48932 4282 48988
rect 4282 48932 4338 48988
rect 4338 48932 4342 48988
rect 4278 48928 4342 48932
rect 4358 48988 4422 48992
rect 4358 48932 4362 48988
rect 4362 48932 4418 48988
rect 4418 48932 4422 48988
rect 4358 48928 4422 48932
rect 4438 48988 4502 48992
rect 4438 48932 4442 48988
rect 4442 48932 4498 48988
rect 4498 48932 4502 48988
rect 4438 48928 4502 48932
rect 34918 48988 34982 48992
rect 34918 48932 34922 48988
rect 34922 48932 34978 48988
rect 34978 48932 34982 48988
rect 34918 48928 34982 48932
rect 34998 48988 35062 48992
rect 34998 48932 35002 48988
rect 35002 48932 35058 48988
rect 35058 48932 35062 48988
rect 34998 48928 35062 48932
rect 35078 48988 35142 48992
rect 35078 48932 35082 48988
rect 35082 48932 35138 48988
rect 35138 48932 35142 48988
rect 35078 48928 35142 48932
rect 35158 48988 35222 48992
rect 35158 48932 35162 48988
rect 35162 48932 35218 48988
rect 35218 48932 35222 48988
rect 35158 48928 35222 48932
rect 19558 48444 19622 48448
rect 19558 48388 19562 48444
rect 19562 48388 19618 48444
rect 19618 48388 19622 48444
rect 19558 48384 19622 48388
rect 19638 48444 19702 48448
rect 19638 48388 19642 48444
rect 19642 48388 19698 48444
rect 19698 48388 19702 48444
rect 19638 48384 19702 48388
rect 19718 48444 19782 48448
rect 19718 48388 19722 48444
rect 19722 48388 19778 48444
rect 19778 48388 19782 48444
rect 19718 48384 19782 48388
rect 19798 48444 19862 48448
rect 19798 48388 19802 48444
rect 19802 48388 19858 48444
rect 19858 48388 19862 48444
rect 19798 48384 19862 48388
rect 50278 48444 50342 48448
rect 50278 48388 50282 48444
rect 50282 48388 50338 48444
rect 50338 48388 50342 48444
rect 50278 48384 50342 48388
rect 50358 48444 50422 48448
rect 50358 48388 50362 48444
rect 50362 48388 50418 48444
rect 50418 48388 50422 48444
rect 50358 48384 50422 48388
rect 50438 48444 50502 48448
rect 50438 48388 50442 48444
rect 50442 48388 50498 48444
rect 50498 48388 50502 48444
rect 50438 48384 50502 48388
rect 50518 48444 50582 48448
rect 50518 48388 50522 48444
rect 50522 48388 50578 48444
rect 50578 48388 50582 48444
rect 50518 48384 50582 48388
rect 4198 47900 4262 47904
rect 4198 47844 4202 47900
rect 4202 47844 4258 47900
rect 4258 47844 4262 47900
rect 4198 47840 4262 47844
rect 4278 47900 4342 47904
rect 4278 47844 4282 47900
rect 4282 47844 4338 47900
rect 4338 47844 4342 47900
rect 4278 47840 4342 47844
rect 4358 47900 4422 47904
rect 4358 47844 4362 47900
rect 4362 47844 4418 47900
rect 4418 47844 4422 47900
rect 4358 47840 4422 47844
rect 4438 47900 4502 47904
rect 4438 47844 4442 47900
rect 4442 47844 4498 47900
rect 4498 47844 4502 47900
rect 4438 47840 4502 47844
rect 34918 47900 34982 47904
rect 34918 47844 34922 47900
rect 34922 47844 34978 47900
rect 34978 47844 34982 47900
rect 34918 47840 34982 47844
rect 34998 47900 35062 47904
rect 34998 47844 35002 47900
rect 35002 47844 35058 47900
rect 35058 47844 35062 47900
rect 34998 47840 35062 47844
rect 35078 47900 35142 47904
rect 35078 47844 35082 47900
rect 35082 47844 35138 47900
rect 35138 47844 35142 47900
rect 35078 47840 35142 47844
rect 35158 47900 35222 47904
rect 35158 47844 35162 47900
rect 35162 47844 35218 47900
rect 35218 47844 35222 47900
rect 35158 47840 35222 47844
rect 19558 47356 19622 47360
rect 19558 47300 19562 47356
rect 19562 47300 19618 47356
rect 19618 47300 19622 47356
rect 19558 47296 19622 47300
rect 19638 47356 19702 47360
rect 19638 47300 19642 47356
rect 19642 47300 19698 47356
rect 19698 47300 19702 47356
rect 19638 47296 19702 47300
rect 19718 47356 19782 47360
rect 19718 47300 19722 47356
rect 19722 47300 19778 47356
rect 19778 47300 19782 47356
rect 19718 47296 19782 47300
rect 19798 47356 19862 47360
rect 19798 47300 19802 47356
rect 19802 47300 19858 47356
rect 19858 47300 19862 47356
rect 19798 47296 19862 47300
rect 50278 47356 50342 47360
rect 50278 47300 50282 47356
rect 50282 47300 50338 47356
rect 50338 47300 50342 47356
rect 50278 47296 50342 47300
rect 50358 47356 50422 47360
rect 50358 47300 50362 47356
rect 50362 47300 50418 47356
rect 50418 47300 50422 47356
rect 50358 47296 50422 47300
rect 50438 47356 50502 47360
rect 50438 47300 50442 47356
rect 50442 47300 50498 47356
rect 50498 47300 50502 47356
rect 50438 47296 50502 47300
rect 50518 47356 50582 47360
rect 50518 47300 50522 47356
rect 50522 47300 50578 47356
rect 50578 47300 50582 47356
rect 50518 47296 50582 47300
rect 4198 46812 4262 46816
rect 4198 46756 4202 46812
rect 4202 46756 4258 46812
rect 4258 46756 4262 46812
rect 4198 46752 4262 46756
rect 4278 46812 4342 46816
rect 4278 46756 4282 46812
rect 4282 46756 4338 46812
rect 4338 46756 4342 46812
rect 4278 46752 4342 46756
rect 4358 46812 4422 46816
rect 4358 46756 4362 46812
rect 4362 46756 4418 46812
rect 4418 46756 4422 46812
rect 4358 46752 4422 46756
rect 4438 46812 4502 46816
rect 4438 46756 4442 46812
rect 4442 46756 4498 46812
rect 4498 46756 4502 46812
rect 4438 46752 4502 46756
rect 34918 46812 34982 46816
rect 34918 46756 34922 46812
rect 34922 46756 34978 46812
rect 34978 46756 34982 46812
rect 34918 46752 34982 46756
rect 34998 46812 35062 46816
rect 34998 46756 35002 46812
rect 35002 46756 35058 46812
rect 35058 46756 35062 46812
rect 34998 46752 35062 46756
rect 35078 46812 35142 46816
rect 35078 46756 35082 46812
rect 35082 46756 35138 46812
rect 35138 46756 35142 46812
rect 35078 46752 35142 46756
rect 35158 46812 35222 46816
rect 35158 46756 35162 46812
rect 35162 46756 35218 46812
rect 35218 46756 35222 46812
rect 35158 46752 35222 46756
rect 19558 46268 19622 46272
rect 19558 46212 19562 46268
rect 19562 46212 19618 46268
rect 19618 46212 19622 46268
rect 19558 46208 19622 46212
rect 19638 46268 19702 46272
rect 19638 46212 19642 46268
rect 19642 46212 19698 46268
rect 19698 46212 19702 46268
rect 19638 46208 19702 46212
rect 19718 46268 19782 46272
rect 19718 46212 19722 46268
rect 19722 46212 19778 46268
rect 19778 46212 19782 46268
rect 19718 46208 19782 46212
rect 19798 46268 19862 46272
rect 19798 46212 19802 46268
rect 19802 46212 19858 46268
rect 19858 46212 19862 46268
rect 19798 46208 19862 46212
rect 50278 46268 50342 46272
rect 50278 46212 50282 46268
rect 50282 46212 50338 46268
rect 50338 46212 50342 46268
rect 50278 46208 50342 46212
rect 50358 46268 50422 46272
rect 50358 46212 50362 46268
rect 50362 46212 50418 46268
rect 50418 46212 50422 46268
rect 50358 46208 50422 46212
rect 50438 46268 50502 46272
rect 50438 46212 50442 46268
rect 50442 46212 50498 46268
rect 50498 46212 50502 46268
rect 50438 46208 50502 46212
rect 50518 46268 50582 46272
rect 50518 46212 50522 46268
rect 50522 46212 50578 46268
rect 50578 46212 50582 46268
rect 50518 46208 50582 46212
rect 4198 45724 4262 45728
rect 4198 45668 4202 45724
rect 4202 45668 4258 45724
rect 4258 45668 4262 45724
rect 4198 45664 4262 45668
rect 4278 45724 4342 45728
rect 4278 45668 4282 45724
rect 4282 45668 4338 45724
rect 4338 45668 4342 45724
rect 4278 45664 4342 45668
rect 4358 45724 4422 45728
rect 4358 45668 4362 45724
rect 4362 45668 4418 45724
rect 4418 45668 4422 45724
rect 4358 45664 4422 45668
rect 4438 45724 4502 45728
rect 4438 45668 4442 45724
rect 4442 45668 4498 45724
rect 4498 45668 4502 45724
rect 4438 45664 4502 45668
rect 34918 45724 34982 45728
rect 34918 45668 34922 45724
rect 34922 45668 34978 45724
rect 34978 45668 34982 45724
rect 34918 45664 34982 45668
rect 34998 45724 35062 45728
rect 34998 45668 35002 45724
rect 35002 45668 35058 45724
rect 35058 45668 35062 45724
rect 34998 45664 35062 45668
rect 35078 45724 35142 45728
rect 35078 45668 35082 45724
rect 35082 45668 35138 45724
rect 35138 45668 35142 45724
rect 35078 45664 35142 45668
rect 35158 45724 35222 45728
rect 35158 45668 35162 45724
rect 35162 45668 35218 45724
rect 35218 45668 35222 45724
rect 35158 45664 35222 45668
rect 19558 45180 19622 45184
rect 19558 45124 19562 45180
rect 19562 45124 19618 45180
rect 19618 45124 19622 45180
rect 19558 45120 19622 45124
rect 19638 45180 19702 45184
rect 19638 45124 19642 45180
rect 19642 45124 19698 45180
rect 19698 45124 19702 45180
rect 19638 45120 19702 45124
rect 19718 45180 19782 45184
rect 19718 45124 19722 45180
rect 19722 45124 19778 45180
rect 19778 45124 19782 45180
rect 19718 45120 19782 45124
rect 19798 45180 19862 45184
rect 19798 45124 19802 45180
rect 19802 45124 19858 45180
rect 19858 45124 19862 45180
rect 19798 45120 19862 45124
rect 50278 45180 50342 45184
rect 50278 45124 50282 45180
rect 50282 45124 50338 45180
rect 50338 45124 50342 45180
rect 50278 45120 50342 45124
rect 50358 45180 50422 45184
rect 50358 45124 50362 45180
rect 50362 45124 50418 45180
rect 50418 45124 50422 45180
rect 50358 45120 50422 45124
rect 50438 45180 50502 45184
rect 50438 45124 50442 45180
rect 50442 45124 50498 45180
rect 50498 45124 50502 45180
rect 50438 45120 50502 45124
rect 50518 45180 50582 45184
rect 50518 45124 50522 45180
rect 50522 45124 50578 45180
rect 50578 45124 50582 45180
rect 50518 45120 50582 45124
rect 4198 44636 4262 44640
rect 4198 44580 4202 44636
rect 4202 44580 4258 44636
rect 4258 44580 4262 44636
rect 4198 44576 4262 44580
rect 4278 44636 4342 44640
rect 4278 44580 4282 44636
rect 4282 44580 4338 44636
rect 4338 44580 4342 44636
rect 4278 44576 4342 44580
rect 4358 44636 4422 44640
rect 4358 44580 4362 44636
rect 4362 44580 4418 44636
rect 4418 44580 4422 44636
rect 4358 44576 4422 44580
rect 4438 44636 4502 44640
rect 4438 44580 4442 44636
rect 4442 44580 4498 44636
rect 4498 44580 4502 44636
rect 4438 44576 4502 44580
rect 34918 44636 34982 44640
rect 34918 44580 34922 44636
rect 34922 44580 34978 44636
rect 34978 44580 34982 44636
rect 34918 44576 34982 44580
rect 34998 44636 35062 44640
rect 34998 44580 35002 44636
rect 35002 44580 35058 44636
rect 35058 44580 35062 44636
rect 34998 44576 35062 44580
rect 35078 44636 35142 44640
rect 35078 44580 35082 44636
rect 35082 44580 35138 44636
rect 35138 44580 35142 44636
rect 35078 44576 35142 44580
rect 35158 44636 35222 44640
rect 35158 44580 35162 44636
rect 35162 44580 35218 44636
rect 35218 44580 35222 44636
rect 35158 44576 35222 44580
rect 38866 44160 38930 44164
rect 38866 44104 38880 44160
rect 38880 44104 38930 44160
rect 38866 44100 38930 44104
rect 19558 44092 19622 44096
rect 19558 44036 19562 44092
rect 19562 44036 19618 44092
rect 19618 44036 19622 44092
rect 19558 44032 19622 44036
rect 19638 44092 19702 44096
rect 19638 44036 19642 44092
rect 19642 44036 19698 44092
rect 19698 44036 19702 44092
rect 19638 44032 19702 44036
rect 19718 44092 19782 44096
rect 19718 44036 19722 44092
rect 19722 44036 19778 44092
rect 19778 44036 19782 44092
rect 19718 44032 19782 44036
rect 19798 44092 19862 44096
rect 19798 44036 19802 44092
rect 19802 44036 19858 44092
rect 19858 44036 19862 44092
rect 19798 44032 19862 44036
rect 50278 44092 50342 44096
rect 50278 44036 50282 44092
rect 50282 44036 50338 44092
rect 50338 44036 50342 44092
rect 50278 44032 50342 44036
rect 50358 44092 50422 44096
rect 50358 44036 50362 44092
rect 50362 44036 50418 44092
rect 50418 44036 50422 44092
rect 50358 44032 50422 44036
rect 50438 44092 50502 44096
rect 50438 44036 50442 44092
rect 50442 44036 50498 44092
rect 50498 44036 50502 44092
rect 50438 44032 50502 44036
rect 50518 44092 50582 44096
rect 50518 44036 50522 44092
rect 50522 44036 50578 44092
rect 50578 44036 50582 44092
rect 50518 44032 50582 44036
rect 4198 43548 4262 43552
rect 4198 43492 4202 43548
rect 4202 43492 4258 43548
rect 4258 43492 4262 43548
rect 4198 43488 4262 43492
rect 4278 43548 4342 43552
rect 4278 43492 4282 43548
rect 4282 43492 4338 43548
rect 4338 43492 4342 43548
rect 4278 43488 4342 43492
rect 4358 43548 4422 43552
rect 4358 43492 4362 43548
rect 4362 43492 4418 43548
rect 4418 43492 4422 43548
rect 4358 43488 4422 43492
rect 4438 43548 4502 43552
rect 4438 43492 4442 43548
rect 4442 43492 4498 43548
rect 4498 43492 4502 43548
rect 4438 43488 4502 43492
rect 34918 43548 34982 43552
rect 34918 43492 34922 43548
rect 34922 43492 34978 43548
rect 34978 43492 34982 43548
rect 34918 43488 34982 43492
rect 34998 43548 35062 43552
rect 34998 43492 35002 43548
rect 35002 43492 35058 43548
rect 35058 43492 35062 43548
rect 34998 43488 35062 43492
rect 35078 43548 35142 43552
rect 35078 43492 35082 43548
rect 35082 43492 35138 43548
rect 35138 43492 35142 43548
rect 35078 43488 35142 43492
rect 35158 43548 35222 43552
rect 35158 43492 35162 43548
rect 35162 43492 35218 43548
rect 35218 43492 35222 43548
rect 35158 43488 35222 43492
rect 19558 43004 19622 43008
rect 19558 42948 19562 43004
rect 19562 42948 19618 43004
rect 19618 42948 19622 43004
rect 19558 42944 19622 42948
rect 19638 43004 19702 43008
rect 19638 42948 19642 43004
rect 19642 42948 19698 43004
rect 19698 42948 19702 43004
rect 19638 42944 19702 42948
rect 19718 43004 19782 43008
rect 19718 42948 19722 43004
rect 19722 42948 19778 43004
rect 19778 42948 19782 43004
rect 19718 42944 19782 42948
rect 19798 43004 19862 43008
rect 19798 42948 19802 43004
rect 19802 42948 19858 43004
rect 19858 42948 19862 43004
rect 19798 42944 19862 42948
rect 50278 43004 50342 43008
rect 50278 42948 50282 43004
rect 50282 42948 50338 43004
rect 50338 42948 50342 43004
rect 50278 42944 50342 42948
rect 50358 43004 50422 43008
rect 50358 42948 50362 43004
rect 50362 42948 50418 43004
rect 50418 42948 50422 43004
rect 50358 42944 50422 42948
rect 50438 43004 50502 43008
rect 50438 42948 50442 43004
rect 50442 42948 50498 43004
rect 50498 42948 50502 43004
rect 50438 42944 50502 42948
rect 50518 43004 50582 43008
rect 50518 42948 50522 43004
rect 50522 42948 50578 43004
rect 50578 42948 50582 43004
rect 50518 42944 50582 42948
rect 4198 42460 4262 42464
rect 4198 42404 4202 42460
rect 4202 42404 4258 42460
rect 4258 42404 4262 42460
rect 4198 42400 4262 42404
rect 4278 42460 4342 42464
rect 4278 42404 4282 42460
rect 4282 42404 4338 42460
rect 4338 42404 4342 42460
rect 4278 42400 4342 42404
rect 4358 42460 4422 42464
rect 4358 42404 4362 42460
rect 4362 42404 4418 42460
rect 4418 42404 4422 42460
rect 4358 42400 4422 42404
rect 4438 42460 4502 42464
rect 4438 42404 4442 42460
rect 4442 42404 4498 42460
rect 4498 42404 4502 42460
rect 4438 42400 4502 42404
rect 34918 42460 34982 42464
rect 34918 42404 34922 42460
rect 34922 42404 34978 42460
rect 34978 42404 34982 42460
rect 34918 42400 34982 42404
rect 34998 42460 35062 42464
rect 34998 42404 35002 42460
rect 35002 42404 35058 42460
rect 35058 42404 35062 42460
rect 34998 42400 35062 42404
rect 35078 42460 35142 42464
rect 35078 42404 35082 42460
rect 35082 42404 35138 42460
rect 35138 42404 35142 42460
rect 35078 42400 35142 42404
rect 35158 42460 35222 42464
rect 35158 42404 35162 42460
rect 35162 42404 35218 42460
rect 35218 42404 35222 42460
rect 35158 42400 35222 42404
rect 19558 41916 19622 41920
rect 19558 41860 19562 41916
rect 19562 41860 19618 41916
rect 19618 41860 19622 41916
rect 19558 41856 19622 41860
rect 19638 41916 19702 41920
rect 19638 41860 19642 41916
rect 19642 41860 19698 41916
rect 19698 41860 19702 41916
rect 19638 41856 19702 41860
rect 19718 41916 19782 41920
rect 19718 41860 19722 41916
rect 19722 41860 19778 41916
rect 19778 41860 19782 41916
rect 19718 41856 19782 41860
rect 19798 41916 19862 41920
rect 19798 41860 19802 41916
rect 19802 41860 19858 41916
rect 19858 41860 19862 41916
rect 19798 41856 19862 41860
rect 50278 41916 50342 41920
rect 50278 41860 50282 41916
rect 50282 41860 50338 41916
rect 50338 41860 50342 41916
rect 50278 41856 50342 41860
rect 50358 41916 50422 41920
rect 50358 41860 50362 41916
rect 50362 41860 50418 41916
rect 50418 41860 50422 41916
rect 50358 41856 50422 41860
rect 50438 41916 50502 41920
rect 50438 41860 50442 41916
rect 50442 41860 50498 41916
rect 50498 41860 50502 41916
rect 50438 41856 50502 41860
rect 50518 41916 50582 41920
rect 50518 41860 50522 41916
rect 50522 41860 50578 41916
rect 50578 41860 50582 41916
rect 50518 41856 50582 41860
rect 4198 41372 4262 41376
rect 4198 41316 4202 41372
rect 4202 41316 4258 41372
rect 4258 41316 4262 41372
rect 4198 41312 4262 41316
rect 4278 41372 4342 41376
rect 4278 41316 4282 41372
rect 4282 41316 4338 41372
rect 4338 41316 4342 41372
rect 4278 41312 4342 41316
rect 4358 41372 4422 41376
rect 4358 41316 4362 41372
rect 4362 41316 4418 41372
rect 4418 41316 4422 41372
rect 4358 41312 4422 41316
rect 4438 41372 4502 41376
rect 4438 41316 4442 41372
rect 4442 41316 4498 41372
rect 4498 41316 4502 41372
rect 4438 41312 4502 41316
rect 34918 41372 34982 41376
rect 34918 41316 34922 41372
rect 34922 41316 34978 41372
rect 34978 41316 34982 41372
rect 34918 41312 34982 41316
rect 34998 41372 35062 41376
rect 34998 41316 35002 41372
rect 35002 41316 35058 41372
rect 35058 41316 35062 41372
rect 34998 41312 35062 41316
rect 35078 41372 35142 41376
rect 35078 41316 35082 41372
rect 35082 41316 35138 41372
rect 35138 41316 35142 41372
rect 35078 41312 35142 41316
rect 35158 41372 35222 41376
rect 35158 41316 35162 41372
rect 35162 41316 35218 41372
rect 35218 41316 35222 41372
rect 35158 41312 35222 41316
rect 19558 40828 19622 40832
rect 19558 40772 19562 40828
rect 19562 40772 19618 40828
rect 19618 40772 19622 40828
rect 19558 40768 19622 40772
rect 19638 40828 19702 40832
rect 19638 40772 19642 40828
rect 19642 40772 19698 40828
rect 19698 40772 19702 40828
rect 19638 40768 19702 40772
rect 19718 40828 19782 40832
rect 19718 40772 19722 40828
rect 19722 40772 19778 40828
rect 19778 40772 19782 40828
rect 19718 40768 19782 40772
rect 19798 40828 19862 40832
rect 19798 40772 19802 40828
rect 19802 40772 19858 40828
rect 19858 40772 19862 40828
rect 19798 40768 19862 40772
rect 50278 40828 50342 40832
rect 50278 40772 50282 40828
rect 50282 40772 50338 40828
rect 50338 40772 50342 40828
rect 50278 40768 50342 40772
rect 50358 40828 50422 40832
rect 50358 40772 50362 40828
rect 50362 40772 50418 40828
rect 50418 40772 50422 40828
rect 50358 40768 50422 40772
rect 50438 40828 50502 40832
rect 50438 40772 50442 40828
rect 50442 40772 50498 40828
rect 50498 40772 50502 40828
rect 50438 40768 50502 40772
rect 50518 40828 50582 40832
rect 50518 40772 50522 40828
rect 50522 40772 50578 40828
rect 50578 40772 50582 40828
rect 50518 40768 50582 40772
rect 4198 40284 4262 40288
rect 4198 40228 4202 40284
rect 4202 40228 4258 40284
rect 4258 40228 4262 40284
rect 4198 40224 4262 40228
rect 4278 40284 4342 40288
rect 4278 40228 4282 40284
rect 4282 40228 4338 40284
rect 4338 40228 4342 40284
rect 4278 40224 4342 40228
rect 4358 40284 4422 40288
rect 4358 40228 4362 40284
rect 4362 40228 4418 40284
rect 4418 40228 4422 40284
rect 4358 40224 4422 40228
rect 4438 40284 4502 40288
rect 4438 40228 4442 40284
rect 4442 40228 4498 40284
rect 4498 40228 4502 40284
rect 4438 40224 4502 40228
rect 34918 40284 34982 40288
rect 34918 40228 34922 40284
rect 34922 40228 34978 40284
rect 34978 40228 34982 40284
rect 34918 40224 34982 40228
rect 34998 40284 35062 40288
rect 34998 40228 35002 40284
rect 35002 40228 35058 40284
rect 35058 40228 35062 40284
rect 34998 40224 35062 40228
rect 35078 40284 35142 40288
rect 35078 40228 35082 40284
rect 35082 40228 35138 40284
rect 35138 40228 35142 40284
rect 35078 40224 35142 40228
rect 35158 40284 35222 40288
rect 35158 40228 35162 40284
rect 35162 40228 35218 40284
rect 35218 40228 35222 40284
rect 35158 40224 35222 40228
rect 19558 39740 19622 39744
rect 19558 39684 19562 39740
rect 19562 39684 19618 39740
rect 19618 39684 19622 39740
rect 19558 39680 19622 39684
rect 19638 39740 19702 39744
rect 19638 39684 19642 39740
rect 19642 39684 19698 39740
rect 19698 39684 19702 39740
rect 19638 39680 19702 39684
rect 19718 39740 19782 39744
rect 19718 39684 19722 39740
rect 19722 39684 19778 39740
rect 19778 39684 19782 39740
rect 19718 39680 19782 39684
rect 19798 39740 19862 39744
rect 19798 39684 19802 39740
rect 19802 39684 19858 39740
rect 19858 39684 19862 39740
rect 19798 39680 19862 39684
rect 50278 39740 50342 39744
rect 50278 39684 50282 39740
rect 50282 39684 50338 39740
rect 50338 39684 50342 39740
rect 50278 39680 50342 39684
rect 50358 39740 50422 39744
rect 50358 39684 50362 39740
rect 50362 39684 50418 39740
rect 50418 39684 50422 39740
rect 50358 39680 50422 39684
rect 50438 39740 50502 39744
rect 50438 39684 50442 39740
rect 50442 39684 50498 39740
rect 50498 39684 50502 39740
rect 50438 39680 50502 39684
rect 50518 39740 50582 39744
rect 50518 39684 50522 39740
rect 50522 39684 50578 39740
rect 50578 39684 50582 39740
rect 50518 39680 50582 39684
rect 4198 39196 4262 39200
rect 4198 39140 4202 39196
rect 4202 39140 4258 39196
rect 4258 39140 4262 39196
rect 4198 39136 4262 39140
rect 4278 39196 4342 39200
rect 4278 39140 4282 39196
rect 4282 39140 4338 39196
rect 4338 39140 4342 39196
rect 4278 39136 4342 39140
rect 4358 39196 4422 39200
rect 4358 39140 4362 39196
rect 4362 39140 4418 39196
rect 4418 39140 4422 39196
rect 4358 39136 4422 39140
rect 4438 39196 4502 39200
rect 4438 39140 4442 39196
rect 4442 39140 4498 39196
rect 4498 39140 4502 39196
rect 4438 39136 4502 39140
rect 34918 39196 34982 39200
rect 34918 39140 34922 39196
rect 34922 39140 34978 39196
rect 34978 39140 34982 39196
rect 34918 39136 34982 39140
rect 34998 39196 35062 39200
rect 34998 39140 35002 39196
rect 35002 39140 35058 39196
rect 35058 39140 35062 39196
rect 34998 39136 35062 39140
rect 35078 39196 35142 39200
rect 35078 39140 35082 39196
rect 35082 39140 35138 39196
rect 35138 39140 35142 39196
rect 35078 39136 35142 39140
rect 35158 39196 35222 39200
rect 35158 39140 35162 39196
rect 35162 39140 35218 39196
rect 35218 39140 35222 39196
rect 35158 39136 35222 39140
rect 19558 38652 19622 38656
rect 19558 38596 19562 38652
rect 19562 38596 19618 38652
rect 19618 38596 19622 38652
rect 19558 38592 19622 38596
rect 19638 38652 19702 38656
rect 19638 38596 19642 38652
rect 19642 38596 19698 38652
rect 19698 38596 19702 38652
rect 19638 38592 19702 38596
rect 19718 38652 19782 38656
rect 19718 38596 19722 38652
rect 19722 38596 19778 38652
rect 19778 38596 19782 38652
rect 19718 38592 19782 38596
rect 19798 38652 19862 38656
rect 19798 38596 19802 38652
rect 19802 38596 19858 38652
rect 19858 38596 19862 38652
rect 19798 38592 19862 38596
rect 50278 38652 50342 38656
rect 50278 38596 50282 38652
rect 50282 38596 50338 38652
rect 50338 38596 50342 38652
rect 50278 38592 50342 38596
rect 50358 38652 50422 38656
rect 50358 38596 50362 38652
rect 50362 38596 50418 38652
rect 50418 38596 50422 38652
rect 50358 38592 50422 38596
rect 50438 38652 50502 38656
rect 50438 38596 50442 38652
rect 50442 38596 50498 38652
rect 50498 38596 50502 38652
rect 50438 38592 50502 38596
rect 50518 38652 50582 38656
rect 50518 38596 50522 38652
rect 50522 38596 50578 38652
rect 50578 38596 50582 38652
rect 50518 38592 50582 38596
rect 4198 38108 4262 38112
rect 4198 38052 4202 38108
rect 4202 38052 4258 38108
rect 4258 38052 4262 38108
rect 4198 38048 4262 38052
rect 4278 38108 4342 38112
rect 4278 38052 4282 38108
rect 4282 38052 4338 38108
rect 4338 38052 4342 38108
rect 4278 38048 4342 38052
rect 4358 38108 4422 38112
rect 4358 38052 4362 38108
rect 4362 38052 4418 38108
rect 4418 38052 4422 38108
rect 4358 38048 4422 38052
rect 4438 38108 4502 38112
rect 4438 38052 4442 38108
rect 4442 38052 4498 38108
rect 4498 38052 4502 38108
rect 4438 38048 4502 38052
rect 34918 38108 34982 38112
rect 34918 38052 34922 38108
rect 34922 38052 34978 38108
rect 34978 38052 34982 38108
rect 34918 38048 34982 38052
rect 34998 38108 35062 38112
rect 34998 38052 35002 38108
rect 35002 38052 35058 38108
rect 35058 38052 35062 38108
rect 34998 38048 35062 38052
rect 35078 38108 35142 38112
rect 35078 38052 35082 38108
rect 35082 38052 35138 38108
rect 35138 38052 35142 38108
rect 35078 38048 35142 38052
rect 35158 38108 35222 38112
rect 35158 38052 35162 38108
rect 35162 38052 35218 38108
rect 35218 38052 35222 38108
rect 35158 38048 35222 38052
rect 19558 37564 19622 37568
rect 19558 37508 19562 37564
rect 19562 37508 19618 37564
rect 19618 37508 19622 37564
rect 19558 37504 19622 37508
rect 19638 37564 19702 37568
rect 19638 37508 19642 37564
rect 19642 37508 19698 37564
rect 19698 37508 19702 37564
rect 19638 37504 19702 37508
rect 19718 37564 19782 37568
rect 19718 37508 19722 37564
rect 19722 37508 19778 37564
rect 19778 37508 19782 37564
rect 19718 37504 19782 37508
rect 19798 37564 19862 37568
rect 19798 37508 19802 37564
rect 19802 37508 19858 37564
rect 19858 37508 19862 37564
rect 19798 37504 19862 37508
rect 50278 37564 50342 37568
rect 50278 37508 50282 37564
rect 50282 37508 50338 37564
rect 50338 37508 50342 37564
rect 50278 37504 50342 37508
rect 50358 37564 50422 37568
rect 50358 37508 50362 37564
rect 50362 37508 50418 37564
rect 50418 37508 50422 37564
rect 50358 37504 50422 37508
rect 50438 37564 50502 37568
rect 50438 37508 50442 37564
rect 50442 37508 50498 37564
rect 50498 37508 50502 37564
rect 50438 37504 50502 37508
rect 50518 37564 50582 37568
rect 50518 37508 50522 37564
rect 50522 37508 50578 37564
rect 50578 37508 50582 37564
rect 50518 37504 50582 37508
rect 4198 37020 4262 37024
rect 4198 36964 4202 37020
rect 4202 36964 4258 37020
rect 4258 36964 4262 37020
rect 4198 36960 4262 36964
rect 4278 37020 4342 37024
rect 4278 36964 4282 37020
rect 4282 36964 4338 37020
rect 4338 36964 4342 37020
rect 4278 36960 4342 36964
rect 4358 37020 4422 37024
rect 4358 36964 4362 37020
rect 4362 36964 4418 37020
rect 4418 36964 4422 37020
rect 4358 36960 4422 36964
rect 4438 37020 4502 37024
rect 4438 36964 4442 37020
rect 4442 36964 4498 37020
rect 4498 36964 4502 37020
rect 4438 36960 4502 36964
rect 34918 37020 34982 37024
rect 34918 36964 34922 37020
rect 34922 36964 34978 37020
rect 34978 36964 34982 37020
rect 34918 36960 34982 36964
rect 34998 37020 35062 37024
rect 34998 36964 35002 37020
rect 35002 36964 35058 37020
rect 35058 36964 35062 37020
rect 34998 36960 35062 36964
rect 35078 37020 35142 37024
rect 35078 36964 35082 37020
rect 35082 36964 35138 37020
rect 35138 36964 35142 37020
rect 35078 36960 35142 36964
rect 35158 37020 35222 37024
rect 35158 36964 35162 37020
rect 35162 36964 35218 37020
rect 35218 36964 35222 37020
rect 35158 36960 35222 36964
rect 19558 36476 19622 36480
rect 19558 36420 19562 36476
rect 19562 36420 19618 36476
rect 19618 36420 19622 36476
rect 19558 36416 19622 36420
rect 19638 36476 19702 36480
rect 19638 36420 19642 36476
rect 19642 36420 19698 36476
rect 19698 36420 19702 36476
rect 19638 36416 19702 36420
rect 19718 36476 19782 36480
rect 19718 36420 19722 36476
rect 19722 36420 19778 36476
rect 19778 36420 19782 36476
rect 19718 36416 19782 36420
rect 19798 36476 19862 36480
rect 19798 36420 19802 36476
rect 19802 36420 19858 36476
rect 19858 36420 19862 36476
rect 19798 36416 19862 36420
rect 50278 36476 50342 36480
rect 50278 36420 50282 36476
rect 50282 36420 50338 36476
rect 50338 36420 50342 36476
rect 50278 36416 50342 36420
rect 50358 36476 50422 36480
rect 50358 36420 50362 36476
rect 50362 36420 50418 36476
rect 50418 36420 50422 36476
rect 50358 36416 50422 36420
rect 50438 36476 50502 36480
rect 50438 36420 50442 36476
rect 50442 36420 50498 36476
rect 50498 36420 50502 36476
rect 50438 36416 50502 36420
rect 50518 36476 50582 36480
rect 50518 36420 50522 36476
rect 50522 36420 50578 36476
rect 50578 36420 50582 36476
rect 50518 36416 50582 36420
rect 4198 35932 4262 35936
rect 4198 35876 4202 35932
rect 4202 35876 4258 35932
rect 4258 35876 4262 35932
rect 4198 35872 4262 35876
rect 4278 35932 4342 35936
rect 4278 35876 4282 35932
rect 4282 35876 4338 35932
rect 4338 35876 4342 35932
rect 4278 35872 4342 35876
rect 4358 35932 4422 35936
rect 4358 35876 4362 35932
rect 4362 35876 4418 35932
rect 4418 35876 4422 35932
rect 4358 35872 4422 35876
rect 4438 35932 4502 35936
rect 4438 35876 4442 35932
rect 4442 35876 4498 35932
rect 4498 35876 4502 35932
rect 4438 35872 4502 35876
rect 34918 35932 34982 35936
rect 34918 35876 34922 35932
rect 34922 35876 34978 35932
rect 34978 35876 34982 35932
rect 34918 35872 34982 35876
rect 34998 35932 35062 35936
rect 34998 35876 35002 35932
rect 35002 35876 35058 35932
rect 35058 35876 35062 35932
rect 34998 35872 35062 35876
rect 35078 35932 35142 35936
rect 35078 35876 35082 35932
rect 35082 35876 35138 35932
rect 35138 35876 35142 35932
rect 35078 35872 35142 35876
rect 35158 35932 35222 35936
rect 35158 35876 35162 35932
rect 35162 35876 35218 35932
rect 35218 35876 35222 35932
rect 35158 35872 35222 35876
rect 19558 35388 19622 35392
rect 19558 35332 19562 35388
rect 19562 35332 19618 35388
rect 19618 35332 19622 35388
rect 19558 35328 19622 35332
rect 19638 35388 19702 35392
rect 19638 35332 19642 35388
rect 19642 35332 19698 35388
rect 19698 35332 19702 35388
rect 19638 35328 19702 35332
rect 19718 35388 19782 35392
rect 19718 35332 19722 35388
rect 19722 35332 19778 35388
rect 19778 35332 19782 35388
rect 19718 35328 19782 35332
rect 19798 35388 19862 35392
rect 19798 35332 19802 35388
rect 19802 35332 19858 35388
rect 19858 35332 19862 35388
rect 19798 35328 19862 35332
rect 50278 35388 50342 35392
rect 50278 35332 50282 35388
rect 50282 35332 50338 35388
rect 50338 35332 50342 35388
rect 50278 35328 50342 35332
rect 50358 35388 50422 35392
rect 50358 35332 50362 35388
rect 50362 35332 50418 35388
rect 50418 35332 50422 35388
rect 50358 35328 50422 35332
rect 50438 35388 50502 35392
rect 50438 35332 50442 35388
rect 50442 35332 50498 35388
rect 50498 35332 50502 35388
rect 50438 35328 50502 35332
rect 50518 35388 50582 35392
rect 50518 35332 50522 35388
rect 50522 35332 50578 35388
rect 50578 35332 50582 35388
rect 50518 35328 50582 35332
rect 4198 34844 4262 34848
rect 4198 34788 4202 34844
rect 4202 34788 4258 34844
rect 4258 34788 4262 34844
rect 4198 34784 4262 34788
rect 4278 34844 4342 34848
rect 4278 34788 4282 34844
rect 4282 34788 4338 34844
rect 4338 34788 4342 34844
rect 4278 34784 4342 34788
rect 4358 34844 4422 34848
rect 4358 34788 4362 34844
rect 4362 34788 4418 34844
rect 4418 34788 4422 34844
rect 4358 34784 4422 34788
rect 4438 34844 4502 34848
rect 4438 34788 4442 34844
rect 4442 34788 4498 34844
rect 4498 34788 4502 34844
rect 4438 34784 4502 34788
rect 34918 34844 34982 34848
rect 34918 34788 34922 34844
rect 34922 34788 34978 34844
rect 34978 34788 34982 34844
rect 34918 34784 34982 34788
rect 34998 34844 35062 34848
rect 34998 34788 35002 34844
rect 35002 34788 35058 34844
rect 35058 34788 35062 34844
rect 34998 34784 35062 34788
rect 35078 34844 35142 34848
rect 35078 34788 35082 34844
rect 35082 34788 35138 34844
rect 35138 34788 35142 34844
rect 35078 34784 35142 34788
rect 35158 34844 35222 34848
rect 35158 34788 35162 34844
rect 35162 34788 35218 34844
rect 35218 34788 35222 34844
rect 35158 34784 35222 34788
rect 19558 34300 19622 34304
rect 19558 34244 19562 34300
rect 19562 34244 19618 34300
rect 19618 34244 19622 34300
rect 19558 34240 19622 34244
rect 19638 34300 19702 34304
rect 19638 34244 19642 34300
rect 19642 34244 19698 34300
rect 19698 34244 19702 34300
rect 19638 34240 19702 34244
rect 19718 34300 19782 34304
rect 19718 34244 19722 34300
rect 19722 34244 19778 34300
rect 19778 34244 19782 34300
rect 19718 34240 19782 34244
rect 19798 34300 19862 34304
rect 19798 34244 19802 34300
rect 19802 34244 19858 34300
rect 19858 34244 19862 34300
rect 19798 34240 19862 34244
rect 50278 34300 50342 34304
rect 50278 34244 50282 34300
rect 50282 34244 50338 34300
rect 50338 34244 50342 34300
rect 50278 34240 50342 34244
rect 50358 34300 50422 34304
rect 50358 34244 50362 34300
rect 50362 34244 50418 34300
rect 50418 34244 50422 34300
rect 50358 34240 50422 34244
rect 50438 34300 50502 34304
rect 50438 34244 50442 34300
rect 50442 34244 50498 34300
rect 50498 34244 50502 34300
rect 50438 34240 50502 34244
rect 50518 34300 50582 34304
rect 50518 34244 50522 34300
rect 50522 34244 50578 34300
rect 50578 34244 50582 34300
rect 50518 34240 50582 34244
rect 4198 33756 4262 33760
rect 4198 33700 4202 33756
rect 4202 33700 4258 33756
rect 4258 33700 4262 33756
rect 4198 33696 4262 33700
rect 4278 33756 4342 33760
rect 4278 33700 4282 33756
rect 4282 33700 4338 33756
rect 4338 33700 4342 33756
rect 4278 33696 4342 33700
rect 4358 33756 4422 33760
rect 4358 33700 4362 33756
rect 4362 33700 4418 33756
rect 4418 33700 4422 33756
rect 4358 33696 4422 33700
rect 4438 33756 4502 33760
rect 4438 33700 4442 33756
rect 4442 33700 4498 33756
rect 4498 33700 4502 33756
rect 4438 33696 4502 33700
rect 34918 33756 34982 33760
rect 34918 33700 34922 33756
rect 34922 33700 34978 33756
rect 34978 33700 34982 33756
rect 34918 33696 34982 33700
rect 34998 33756 35062 33760
rect 34998 33700 35002 33756
rect 35002 33700 35058 33756
rect 35058 33700 35062 33756
rect 34998 33696 35062 33700
rect 35078 33756 35142 33760
rect 35078 33700 35082 33756
rect 35082 33700 35138 33756
rect 35138 33700 35142 33756
rect 35078 33696 35142 33700
rect 35158 33756 35222 33760
rect 35158 33700 35162 33756
rect 35162 33700 35218 33756
rect 35218 33700 35222 33756
rect 35158 33696 35222 33700
rect 19558 33212 19622 33216
rect 19558 33156 19562 33212
rect 19562 33156 19618 33212
rect 19618 33156 19622 33212
rect 19558 33152 19622 33156
rect 19638 33212 19702 33216
rect 19638 33156 19642 33212
rect 19642 33156 19698 33212
rect 19698 33156 19702 33212
rect 19638 33152 19702 33156
rect 19718 33212 19782 33216
rect 19718 33156 19722 33212
rect 19722 33156 19778 33212
rect 19778 33156 19782 33212
rect 19718 33152 19782 33156
rect 19798 33212 19862 33216
rect 19798 33156 19802 33212
rect 19802 33156 19858 33212
rect 19858 33156 19862 33212
rect 19798 33152 19862 33156
rect 50278 33212 50342 33216
rect 50278 33156 50282 33212
rect 50282 33156 50338 33212
rect 50338 33156 50342 33212
rect 50278 33152 50342 33156
rect 50358 33212 50422 33216
rect 50358 33156 50362 33212
rect 50362 33156 50418 33212
rect 50418 33156 50422 33212
rect 50358 33152 50422 33156
rect 50438 33212 50502 33216
rect 50438 33156 50442 33212
rect 50442 33156 50498 33212
rect 50498 33156 50502 33212
rect 50438 33152 50502 33156
rect 50518 33212 50582 33216
rect 50518 33156 50522 33212
rect 50522 33156 50578 33212
rect 50578 33156 50582 33212
rect 50518 33152 50582 33156
rect 4198 32668 4262 32672
rect 4198 32612 4202 32668
rect 4202 32612 4258 32668
rect 4258 32612 4262 32668
rect 4198 32608 4262 32612
rect 4278 32668 4342 32672
rect 4278 32612 4282 32668
rect 4282 32612 4338 32668
rect 4338 32612 4342 32668
rect 4278 32608 4342 32612
rect 4358 32668 4422 32672
rect 4358 32612 4362 32668
rect 4362 32612 4418 32668
rect 4418 32612 4422 32668
rect 4358 32608 4422 32612
rect 4438 32668 4502 32672
rect 4438 32612 4442 32668
rect 4442 32612 4498 32668
rect 4498 32612 4502 32668
rect 4438 32608 4502 32612
rect 34918 32668 34982 32672
rect 34918 32612 34922 32668
rect 34922 32612 34978 32668
rect 34978 32612 34982 32668
rect 34918 32608 34982 32612
rect 34998 32668 35062 32672
rect 34998 32612 35002 32668
rect 35002 32612 35058 32668
rect 35058 32612 35062 32668
rect 34998 32608 35062 32612
rect 35078 32668 35142 32672
rect 35078 32612 35082 32668
rect 35082 32612 35138 32668
rect 35138 32612 35142 32668
rect 35078 32608 35142 32612
rect 35158 32668 35222 32672
rect 35158 32612 35162 32668
rect 35162 32612 35218 32668
rect 35218 32612 35222 32668
rect 35158 32608 35222 32612
rect 19558 32124 19622 32128
rect 19558 32068 19562 32124
rect 19562 32068 19618 32124
rect 19618 32068 19622 32124
rect 19558 32064 19622 32068
rect 19638 32124 19702 32128
rect 19638 32068 19642 32124
rect 19642 32068 19698 32124
rect 19698 32068 19702 32124
rect 19638 32064 19702 32068
rect 19718 32124 19782 32128
rect 19718 32068 19722 32124
rect 19722 32068 19778 32124
rect 19778 32068 19782 32124
rect 19718 32064 19782 32068
rect 19798 32124 19862 32128
rect 19798 32068 19802 32124
rect 19802 32068 19858 32124
rect 19858 32068 19862 32124
rect 19798 32064 19862 32068
rect 50278 32124 50342 32128
rect 50278 32068 50282 32124
rect 50282 32068 50338 32124
rect 50338 32068 50342 32124
rect 50278 32064 50342 32068
rect 50358 32124 50422 32128
rect 50358 32068 50362 32124
rect 50362 32068 50418 32124
rect 50418 32068 50422 32124
rect 50358 32064 50422 32068
rect 50438 32124 50502 32128
rect 50438 32068 50442 32124
rect 50442 32068 50498 32124
rect 50498 32068 50502 32124
rect 50438 32064 50502 32068
rect 50518 32124 50582 32128
rect 50518 32068 50522 32124
rect 50522 32068 50578 32124
rect 50578 32068 50582 32124
rect 50518 32064 50582 32068
rect 4198 31580 4262 31584
rect 4198 31524 4202 31580
rect 4202 31524 4258 31580
rect 4258 31524 4262 31580
rect 4198 31520 4262 31524
rect 4278 31580 4342 31584
rect 4278 31524 4282 31580
rect 4282 31524 4338 31580
rect 4338 31524 4342 31580
rect 4278 31520 4342 31524
rect 4358 31580 4422 31584
rect 4358 31524 4362 31580
rect 4362 31524 4418 31580
rect 4418 31524 4422 31580
rect 4358 31520 4422 31524
rect 4438 31580 4502 31584
rect 4438 31524 4442 31580
rect 4442 31524 4498 31580
rect 4498 31524 4502 31580
rect 4438 31520 4502 31524
rect 34918 31580 34982 31584
rect 34918 31524 34922 31580
rect 34922 31524 34978 31580
rect 34978 31524 34982 31580
rect 34918 31520 34982 31524
rect 34998 31580 35062 31584
rect 34998 31524 35002 31580
rect 35002 31524 35058 31580
rect 35058 31524 35062 31580
rect 34998 31520 35062 31524
rect 35078 31580 35142 31584
rect 35078 31524 35082 31580
rect 35082 31524 35138 31580
rect 35138 31524 35142 31580
rect 35078 31520 35142 31524
rect 35158 31580 35222 31584
rect 35158 31524 35162 31580
rect 35162 31524 35218 31580
rect 35218 31524 35222 31580
rect 35158 31520 35222 31524
rect 19558 31036 19622 31040
rect 19558 30980 19562 31036
rect 19562 30980 19618 31036
rect 19618 30980 19622 31036
rect 19558 30976 19622 30980
rect 19638 31036 19702 31040
rect 19638 30980 19642 31036
rect 19642 30980 19698 31036
rect 19698 30980 19702 31036
rect 19638 30976 19702 30980
rect 19718 31036 19782 31040
rect 19718 30980 19722 31036
rect 19722 30980 19778 31036
rect 19778 30980 19782 31036
rect 19718 30976 19782 30980
rect 19798 31036 19862 31040
rect 19798 30980 19802 31036
rect 19802 30980 19858 31036
rect 19858 30980 19862 31036
rect 19798 30976 19862 30980
rect 50278 31036 50342 31040
rect 50278 30980 50282 31036
rect 50282 30980 50338 31036
rect 50338 30980 50342 31036
rect 50278 30976 50342 30980
rect 50358 31036 50422 31040
rect 50358 30980 50362 31036
rect 50362 30980 50418 31036
rect 50418 30980 50422 31036
rect 50358 30976 50422 30980
rect 50438 31036 50502 31040
rect 50438 30980 50442 31036
rect 50442 30980 50498 31036
rect 50498 30980 50502 31036
rect 50438 30976 50502 30980
rect 50518 31036 50582 31040
rect 50518 30980 50522 31036
rect 50522 30980 50578 31036
rect 50578 30980 50582 31036
rect 50518 30976 50582 30980
rect 4198 30492 4262 30496
rect 4198 30436 4202 30492
rect 4202 30436 4258 30492
rect 4258 30436 4262 30492
rect 4198 30432 4262 30436
rect 4278 30492 4342 30496
rect 4278 30436 4282 30492
rect 4282 30436 4338 30492
rect 4338 30436 4342 30492
rect 4278 30432 4342 30436
rect 4358 30492 4422 30496
rect 4358 30436 4362 30492
rect 4362 30436 4418 30492
rect 4418 30436 4422 30492
rect 4358 30432 4422 30436
rect 4438 30492 4502 30496
rect 4438 30436 4442 30492
rect 4442 30436 4498 30492
rect 4498 30436 4502 30492
rect 4438 30432 4502 30436
rect 34918 30492 34982 30496
rect 34918 30436 34922 30492
rect 34922 30436 34978 30492
rect 34978 30436 34982 30492
rect 34918 30432 34982 30436
rect 34998 30492 35062 30496
rect 34998 30436 35002 30492
rect 35002 30436 35058 30492
rect 35058 30436 35062 30492
rect 34998 30432 35062 30436
rect 35078 30492 35142 30496
rect 35078 30436 35082 30492
rect 35082 30436 35138 30492
rect 35138 30436 35142 30492
rect 35078 30432 35142 30436
rect 35158 30492 35222 30496
rect 35158 30436 35162 30492
rect 35162 30436 35218 30492
rect 35218 30436 35222 30492
rect 35158 30432 35222 30436
rect 19558 29948 19622 29952
rect 19558 29892 19562 29948
rect 19562 29892 19618 29948
rect 19618 29892 19622 29948
rect 19558 29888 19622 29892
rect 19638 29948 19702 29952
rect 19638 29892 19642 29948
rect 19642 29892 19698 29948
rect 19698 29892 19702 29948
rect 19638 29888 19702 29892
rect 19718 29948 19782 29952
rect 19718 29892 19722 29948
rect 19722 29892 19778 29948
rect 19778 29892 19782 29948
rect 19718 29888 19782 29892
rect 19798 29948 19862 29952
rect 19798 29892 19802 29948
rect 19802 29892 19858 29948
rect 19858 29892 19862 29948
rect 19798 29888 19862 29892
rect 50278 29948 50342 29952
rect 50278 29892 50282 29948
rect 50282 29892 50338 29948
rect 50338 29892 50342 29948
rect 50278 29888 50342 29892
rect 50358 29948 50422 29952
rect 50358 29892 50362 29948
rect 50362 29892 50418 29948
rect 50418 29892 50422 29948
rect 50358 29888 50422 29892
rect 50438 29948 50502 29952
rect 50438 29892 50442 29948
rect 50442 29892 50498 29948
rect 50498 29892 50502 29948
rect 50438 29888 50502 29892
rect 50518 29948 50582 29952
rect 50518 29892 50522 29948
rect 50522 29892 50578 29948
rect 50578 29892 50582 29948
rect 50518 29888 50582 29892
rect 4198 29404 4262 29408
rect 4198 29348 4202 29404
rect 4202 29348 4258 29404
rect 4258 29348 4262 29404
rect 4198 29344 4262 29348
rect 4278 29404 4342 29408
rect 4278 29348 4282 29404
rect 4282 29348 4338 29404
rect 4338 29348 4342 29404
rect 4278 29344 4342 29348
rect 4358 29404 4422 29408
rect 4358 29348 4362 29404
rect 4362 29348 4418 29404
rect 4418 29348 4422 29404
rect 4358 29344 4422 29348
rect 4438 29404 4502 29408
rect 4438 29348 4442 29404
rect 4442 29348 4498 29404
rect 4498 29348 4502 29404
rect 4438 29344 4502 29348
rect 34918 29404 34982 29408
rect 34918 29348 34922 29404
rect 34922 29348 34978 29404
rect 34978 29348 34982 29404
rect 34918 29344 34982 29348
rect 34998 29404 35062 29408
rect 34998 29348 35002 29404
rect 35002 29348 35058 29404
rect 35058 29348 35062 29404
rect 34998 29344 35062 29348
rect 35078 29404 35142 29408
rect 35078 29348 35082 29404
rect 35082 29348 35138 29404
rect 35138 29348 35142 29404
rect 35078 29344 35142 29348
rect 35158 29404 35222 29408
rect 35158 29348 35162 29404
rect 35162 29348 35218 29404
rect 35218 29348 35222 29404
rect 35158 29344 35222 29348
rect 19558 28860 19622 28864
rect 19558 28804 19562 28860
rect 19562 28804 19618 28860
rect 19618 28804 19622 28860
rect 19558 28800 19622 28804
rect 19638 28860 19702 28864
rect 19638 28804 19642 28860
rect 19642 28804 19698 28860
rect 19698 28804 19702 28860
rect 19638 28800 19702 28804
rect 19718 28860 19782 28864
rect 19718 28804 19722 28860
rect 19722 28804 19778 28860
rect 19778 28804 19782 28860
rect 19718 28800 19782 28804
rect 19798 28860 19862 28864
rect 19798 28804 19802 28860
rect 19802 28804 19858 28860
rect 19858 28804 19862 28860
rect 19798 28800 19862 28804
rect 50278 28860 50342 28864
rect 50278 28804 50282 28860
rect 50282 28804 50338 28860
rect 50338 28804 50342 28860
rect 50278 28800 50342 28804
rect 50358 28860 50422 28864
rect 50358 28804 50362 28860
rect 50362 28804 50418 28860
rect 50418 28804 50422 28860
rect 50358 28800 50422 28804
rect 50438 28860 50502 28864
rect 50438 28804 50442 28860
rect 50442 28804 50498 28860
rect 50498 28804 50502 28860
rect 50438 28800 50502 28804
rect 50518 28860 50582 28864
rect 50518 28804 50522 28860
rect 50522 28804 50578 28860
rect 50578 28804 50582 28860
rect 50518 28800 50582 28804
rect 4198 28316 4262 28320
rect 4198 28260 4202 28316
rect 4202 28260 4258 28316
rect 4258 28260 4262 28316
rect 4198 28256 4262 28260
rect 4278 28316 4342 28320
rect 4278 28260 4282 28316
rect 4282 28260 4338 28316
rect 4338 28260 4342 28316
rect 4278 28256 4342 28260
rect 4358 28316 4422 28320
rect 4358 28260 4362 28316
rect 4362 28260 4418 28316
rect 4418 28260 4422 28316
rect 4358 28256 4422 28260
rect 4438 28316 4502 28320
rect 4438 28260 4442 28316
rect 4442 28260 4498 28316
rect 4498 28260 4502 28316
rect 4438 28256 4502 28260
rect 34918 28316 34982 28320
rect 34918 28260 34922 28316
rect 34922 28260 34978 28316
rect 34978 28260 34982 28316
rect 34918 28256 34982 28260
rect 34998 28316 35062 28320
rect 34998 28260 35002 28316
rect 35002 28260 35058 28316
rect 35058 28260 35062 28316
rect 34998 28256 35062 28260
rect 35078 28316 35142 28320
rect 35078 28260 35082 28316
rect 35082 28260 35138 28316
rect 35138 28260 35142 28316
rect 35078 28256 35142 28260
rect 35158 28316 35222 28320
rect 35158 28260 35162 28316
rect 35162 28260 35218 28316
rect 35218 28260 35222 28316
rect 35158 28256 35222 28260
rect 19558 27772 19622 27776
rect 19558 27716 19562 27772
rect 19562 27716 19618 27772
rect 19618 27716 19622 27772
rect 19558 27712 19622 27716
rect 19638 27772 19702 27776
rect 19638 27716 19642 27772
rect 19642 27716 19698 27772
rect 19698 27716 19702 27772
rect 19638 27712 19702 27716
rect 19718 27772 19782 27776
rect 19718 27716 19722 27772
rect 19722 27716 19778 27772
rect 19778 27716 19782 27772
rect 19718 27712 19782 27716
rect 19798 27772 19862 27776
rect 19798 27716 19802 27772
rect 19802 27716 19858 27772
rect 19858 27716 19862 27772
rect 19798 27712 19862 27716
rect 50278 27772 50342 27776
rect 50278 27716 50282 27772
rect 50282 27716 50338 27772
rect 50338 27716 50342 27772
rect 50278 27712 50342 27716
rect 50358 27772 50422 27776
rect 50358 27716 50362 27772
rect 50362 27716 50418 27772
rect 50418 27716 50422 27772
rect 50358 27712 50422 27716
rect 50438 27772 50502 27776
rect 50438 27716 50442 27772
rect 50442 27716 50498 27772
rect 50498 27716 50502 27772
rect 50438 27712 50502 27716
rect 50518 27772 50582 27776
rect 50518 27716 50522 27772
rect 50522 27716 50578 27772
rect 50578 27716 50582 27772
rect 50518 27712 50582 27716
rect 4198 27228 4262 27232
rect 4198 27172 4202 27228
rect 4202 27172 4258 27228
rect 4258 27172 4262 27228
rect 4198 27168 4262 27172
rect 4278 27228 4342 27232
rect 4278 27172 4282 27228
rect 4282 27172 4338 27228
rect 4338 27172 4342 27228
rect 4278 27168 4342 27172
rect 4358 27228 4422 27232
rect 4358 27172 4362 27228
rect 4362 27172 4418 27228
rect 4418 27172 4422 27228
rect 4358 27168 4422 27172
rect 4438 27228 4502 27232
rect 4438 27172 4442 27228
rect 4442 27172 4498 27228
rect 4498 27172 4502 27228
rect 4438 27168 4502 27172
rect 34918 27228 34982 27232
rect 34918 27172 34922 27228
rect 34922 27172 34978 27228
rect 34978 27172 34982 27228
rect 34918 27168 34982 27172
rect 34998 27228 35062 27232
rect 34998 27172 35002 27228
rect 35002 27172 35058 27228
rect 35058 27172 35062 27228
rect 34998 27168 35062 27172
rect 35078 27228 35142 27232
rect 35078 27172 35082 27228
rect 35082 27172 35138 27228
rect 35138 27172 35142 27228
rect 35078 27168 35142 27172
rect 35158 27228 35222 27232
rect 35158 27172 35162 27228
rect 35162 27172 35218 27228
rect 35218 27172 35222 27228
rect 35158 27168 35222 27172
rect 19558 26684 19622 26688
rect 19558 26628 19562 26684
rect 19562 26628 19618 26684
rect 19618 26628 19622 26684
rect 19558 26624 19622 26628
rect 19638 26684 19702 26688
rect 19638 26628 19642 26684
rect 19642 26628 19698 26684
rect 19698 26628 19702 26684
rect 19638 26624 19702 26628
rect 19718 26684 19782 26688
rect 19718 26628 19722 26684
rect 19722 26628 19778 26684
rect 19778 26628 19782 26684
rect 19718 26624 19782 26628
rect 19798 26684 19862 26688
rect 19798 26628 19802 26684
rect 19802 26628 19858 26684
rect 19858 26628 19862 26684
rect 19798 26624 19862 26628
rect 50278 26684 50342 26688
rect 50278 26628 50282 26684
rect 50282 26628 50338 26684
rect 50338 26628 50342 26684
rect 50278 26624 50342 26628
rect 50358 26684 50422 26688
rect 50358 26628 50362 26684
rect 50362 26628 50418 26684
rect 50418 26628 50422 26684
rect 50358 26624 50422 26628
rect 50438 26684 50502 26688
rect 50438 26628 50442 26684
rect 50442 26628 50498 26684
rect 50498 26628 50502 26684
rect 50438 26624 50502 26628
rect 50518 26684 50582 26688
rect 50518 26628 50522 26684
rect 50522 26628 50578 26684
rect 50578 26628 50582 26684
rect 50518 26624 50582 26628
rect 38866 26284 38930 26348
rect 4198 26140 4262 26144
rect 4198 26084 4202 26140
rect 4202 26084 4258 26140
rect 4258 26084 4262 26140
rect 4198 26080 4262 26084
rect 4278 26140 4342 26144
rect 4278 26084 4282 26140
rect 4282 26084 4338 26140
rect 4338 26084 4342 26140
rect 4278 26080 4342 26084
rect 4358 26140 4422 26144
rect 4358 26084 4362 26140
rect 4362 26084 4418 26140
rect 4418 26084 4422 26140
rect 4358 26080 4422 26084
rect 4438 26140 4502 26144
rect 4438 26084 4442 26140
rect 4442 26084 4498 26140
rect 4498 26084 4502 26140
rect 4438 26080 4502 26084
rect 34918 26140 34982 26144
rect 34918 26084 34922 26140
rect 34922 26084 34978 26140
rect 34978 26084 34982 26140
rect 34918 26080 34982 26084
rect 34998 26140 35062 26144
rect 34998 26084 35002 26140
rect 35002 26084 35058 26140
rect 35058 26084 35062 26140
rect 34998 26080 35062 26084
rect 35078 26140 35142 26144
rect 35078 26084 35082 26140
rect 35082 26084 35138 26140
rect 35138 26084 35142 26140
rect 35078 26080 35142 26084
rect 35158 26140 35222 26144
rect 35158 26084 35162 26140
rect 35162 26084 35218 26140
rect 35218 26084 35222 26140
rect 35158 26080 35222 26084
rect 19558 25596 19622 25600
rect 19558 25540 19562 25596
rect 19562 25540 19618 25596
rect 19618 25540 19622 25596
rect 19558 25536 19622 25540
rect 19638 25596 19702 25600
rect 19638 25540 19642 25596
rect 19642 25540 19698 25596
rect 19698 25540 19702 25596
rect 19638 25536 19702 25540
rect 19718 25596 19782 25600
rect 19718 25540 19722 25596
rect 19722 25540 19778 25596
rect 19778 25540 19782 25596
rect 19718 25536 19782 25540
rect 19798 25596 19862 25600
rect 19798 25540 19802 25596
rect 19802 25540 19858 25596
rect 19858 25540 19862 25596
rect 19798 25536 19862 25540
rect 50278 25596 50342 25600
rect 50278 25540 50282 25596
rect 50282 25540 50338 25596
rect 50338 25540 50342 25596
rect 50278 25536 50342 25540
rect 50358 25596 50422 25600
rect 50358 25540 50362 25596
rect 50362 25540 50418 25596
rect 50418 25540 50422 25596
rect 50358 25536 50422 25540
rect 50438 25596 50502 25600
rect 50438 25540 50442 25596
rect 50442 25540 50498 25596
rect 50498 25540 50502 25596
rect 50438 25536 50502 25540
rect 50518 25596 50582 25600
rect 50518 25540 50522 25596
rect 50522 25540 50578 25596
rect 50578 25540 50582 25596
rect 50518 25536 50582 25540
rect 4198 25052 4262 25056
rect 4198 24996 4202 25052
rect 4202 24996 4258 25052
rect 4258 24996 4262 25052
rect 4198 24992 4262 24996
rect 4278 25052 4342 25056
rect 4278 24996 4282 25052
rect 4282 24996 4338 25052
rect 4338 24996 4342 25052
rect 4278 24992 4342 24996
rect 4358 25052 4422 25056
rect 4358 24996 4362 25052
rect 4362 24996 4418 25052
rect 4418 24996 4422 25052
rect 4358 24992 4422 24996
rect 4438 25052 4502 25056
rect 4438 24996 4442 25052
rect 4442 24996 4498 25052
rect 4498 24996 4502 25052
rect 4438 24992 4502 24996
rect 34918 25052 34982 25056
rect 34918 24996 34922 25052
rect 34922 24996 34978 25052
rect 34978 24996 34982 25052
rect 34918 24992 34982 24996
rect 34998 25052 35062 25056
rect 34998 24996 35002 25052
rect 35002 24996 35058 25052
rect 35058 24996 35062 25052
rect 34998 24992 35062 24996
rect 35078 25052 35142 25056
rect 35078 24996 35082 25052
rect 35082 24996 35138 25052
rect 35138 24996 35142 25052
rect 35078 24992 35142 24996
rect 35158 25052 35222 25056
rect 35158 24996 35162 25052
rect 35162 24996 35218 25052
rect 35218 24996 35222 25052
rect 35158 24992 35222 24996
rect 19558 24508 19622 24512
rect 19558 24452 19562 24508
rect 19562 24452 19618 24508
rect 19618 24452 19622 24508
rect 19558 24448 19622 24452
rect 19638 24508 19702 24512
rect 19638 24452 19642 24508
rect 19642 24452 19698 24508
rect 19698 24452 19702 24508
rect 19638 24448 19702 24452
rect 19718 24508 19782 24512
rect 19718 24452 19722 24508
rect 19722 24452 19778 24508
rect 19778 24452 19782 24508
rect 19718 24448 19782 24452
rect 19798 24508 19862 24512
rect 19798 24452 19802 24508
rect 19802 24452 19858 24508
rect 19858 24452 19862 24508
rect 19798 24448 19862 24452
rect 50278 24508 50342 24512
rect 50278 24452 50282 24508
rect 50282 24452 50338 24508
rect 50338 24452 50342 24508
rect 50278 24448 50342 24452
rect 50358 24508 50422 24512
rect 50358 24452 50362 24508
rect 50362 24452 50418 24508
rect 50418 24452 50422 24508
rect 50358 24448 50422 24452
rect 50438 24508 50502 24512
rect 50438 24452 50442 24508
rect 50442 24452 50498 24508
rect 50498 24452 50502 24508
rect 50438 24448 50502 24452
rect 50518 24508 50582 24512
rect 50518 24452 50522 24508
rect 50522 24452 50578 24508
rect 50578 24452 50582 24508
rect 50518 24448 50582 24452
rect 4198 23964 4262 23968
rect 4198 23908 4202 23964
rect 4202 23908 4258 23964
rect 4258 23908 4262 23964
rect 4198 23904 4262 23908
rect 4278 23964 4342 23968
rect 4278 23908 4282 23964
rect 4282 23908 4338 23964
rect 4338 23908 4342 23964
rect 4278 23904 4342 23908
rect 4358 23964 4422 23968
rect 4358 23908 4362 23964
rect 4362 23908 4418 23964
rect 4418 23908 4422 23964
rect 4358 23904 4422 23908
rect 4438 23964 4502 23968
rect 4438 23908 4442 23964
rect 4442 23908 4498 23964
rect 4498 23908 4502 23964
rect 4438 23904 4502 23908
rect 34918 23964 34982 23968
rect 34918 23908 34922 23964
rect 34922 23908 34978 23964
rect 34978 23908 34982 23964
rect 34918 23904 34982 23908
rect 34998 23964 35062 23968
rect 34998 23908 35002 23964
rect 35002 23908 35058 23964
rect 35058 23908 35062 23964
rect 34998 23904 35062 23908
rect 35078 23964 35142 23968
rect 35078 23908 35082 23964
rect 35082 23908 35138 23964
rect 35138 23908 35142 23964
rect 35078 23904 35142 23908
rect 35158 23964 35222 23968
rect 35158 23908 35162 23964
rect 35162 23908 35218 23964
rect 35218 23908 35222 23964
rect 35158 23904 35222 23908
rect 19558 23420 19622 23424
rect 19558 23364 19562 23420
rect 19562 23364 19618 23420
rect 19618 23364 19622 23420
rect 19558 23360 19622 23364
rect 19638 23420 19702 23424
rect 19638 23364 19642 23420
rect 19642 23364 19698 23420
rect 19698 23364 19702 23420
rect 19638 23360 19702 23364
rect 19718 23420 19782 23424
rect 19718 23364 19722 23420
rect 19722 23364 19778 23420
rect 19778 23364 19782 23420
rect 19718 23360 19782 23364
rect 19798 23420 19862 23424
rect 19798 23364 19802 23420
rect 19802 23364 19858 23420
rect 19858 23364 19862 23420
rect 19798 23360 19862 23364
rect 50278 23420 50342 23424
rect 50278 23364 50282 23420
rect 50282 23364 50338 23420
rect 50338 23364 50342 23420
rect 50278 23360 50342 23364
rect 50358 23420 50422 23424
rect 50358 23364 50362 23420
rect 50362 23364 50418 23420
rect 50418 23364 50422 23420
rect 50358 23360 50422 23364
rect 50438 23420 50502 23424
rect 50438 23364 50442 23420
rect 50442 23364 50498 23420
rect 50498 23364 50502 23420
rect 50438 23360 50502 23364
rect 50518 23420 50582 23424
rect 50518 23364 50522 23420
rect 50522 23364 50578 23420
rect 50578 23364 50582 23420
rect 50518 23360 50582 23364
rect 23410 23292 23474 23356
rect 4198 22876 4262 22880
rect 4198 22820 4202 22876
rect 4202 22820 4258 22876
rect 4258 22820 4262 22876
rect 4198 22816 4262 22820
rect 4278 22876 4342 22880
rect 4278 22820 4282 22876
rect 4282 22820 4338 22876
rect 4338 22820 4342 22876
rect 4278 22816 4342 22820
rect 4358 22876 4422 22880
rect 4358 22820 4362 22876
rect 4362 22820 4418 22876
rect 4418 22820 4422 22876
rect 4358 22816 4422 22820
rect 4438 22876 4502 22880
rect 4438 22820 4442 22876
rect 4442 22820 4498 22876
rect 4498 22820 4502 22876
rect 4438 22816 4502 22820
rect 34918 22876 34982 22880
rect 34918 22820 34922 22876
rect 34922 22820 34978 22876
rect 34978 22820 34982 22876
rect 34918 22816 34982 22820
rect 34998 22876 35062 22880
rect 34998 22820 35002 22876
rect 35002 22820 35058 22876
rect 35058 22820 35062 22876
rect 34998 22816 35062 22820
rect 35078 22876 35142 22880
rect 35078 22820 35082 22876
rect 35082 22820 35138 22876
rect 35138 22820 35142 22876
rect 35078 22816 35142 22820
rect 35158 22876 35222 22880
rect 35158 22820 35162 22876
rect 35162 22820 35218 22876
rect 35218 22820 35222 22876
rect 35158 22816 35222 22820
rect 19558 22332 19622 22336
rect 19558 22276 19562 22332
rect 19562 22276 19618 22332
rect 19618 22276 19622 22332
rect 19558 22272 19622 22276
rect 19638 22332 19702 22336
rect 19638 22276 19642 22332
rect 19642 22276 19698 22332
rect 19698 22276 19702 22332
rect 19638 22272 19702 22276
rect 19718 22332 19782 22336
rect 19718 22276 19722 22332
rect 19722 22276 19778 22332
rect 19778 22276 19782 22332
rect 19718 22272 19782 22276
rect 19798 22332 19862 22336
rect 19798 22276 19802 22332
rect 19802 22276 19858 22332
rect 19858 22276 19862 22332
rect 19798 22272 19862 22276
rect 50278 22332 50342 22336
rect 50278 22276 50282 22332
rect 50282 22276 50338 22332
rect 50338 22276 50342 22332
rect 50278 22272 50342 22276
rect 50358 22332 50422 22336
rect 50358 22276 50362 22332
rect 50362 22276 50418 22332
rect 50418 22276 50422 22332
rect 50358 22272 50422 22276
rect 50438 22332 50502 22336
rect 50438 22276 50442 22332
rect 50442 22276 50498 22332
rect 50498 22276 50502 22332
rect 50438 22272 50502 22276
rect 50518 22332 50582 22336
rect 50518 22276 50522 22332
rect 50522 22276 50578 22332
rect 50578 22276 50582 22332
rect 50518 22272 50582 22276
rect 4198 21788 4262 21792
rect 4198 21732 4202 21788
rect 4202 21732 4258 21788
rect 4258 21732 4262 21788
rect 4198 21728 4262 21732
rect 4278 21788 4342 21792
rect 4278 21732 4282 21788
rect 4282 21732 4338 21788
rect 4338 21732 4342 21788
rect 4278 21728 4342 21732
rect 4358 21788 4422 21792
rect 4358 21732 4362 21788
rect 4362 21732 4418 21788
rect 4418 21732 4422 21788
rect 4358 21728 4422 21732
rect 4438 21788 4502 21792
rect 4438 21732 4442 21788
rect 4442 21732 4498 21788
rect 4498 21732 4502 21788
rect 4438 21728 4502 21732
rect 34918 21788 34982 21792
rect 34918 21732 34922 21788
rect 34922 21732 34978 21788
rect 34978 21732 34982 21788
rect 34918 21728 34982 21732
rect 34998 21788 35062 21792
rect 34998 21732 35002 21788
rect 35002 21732 35058 21788
rect 35058 21732 35062 21788
rect 34998 21728 35062 21732
rect 35078 21788 35142 21792
rect 35078 21732 35082 21788
rect 35082 21732 35138 21788
rect 35138 21732 35142 21788
rect 35078 21728 35142 21732
rect 35158 21788 35222 21792
rect 35158 21732 35162 21788
rect 35162 21732 35218 21788
rect 35218 21732 35222 21788
rect 35158 21728 35222 21732
rect 19558 21244 19622 21248
rect 19558 21188 19562 21244
rect 19562 21188 19618 21244
rect 19618 21188 19622 21244
rect 19558 21184 19622 21188
rect 19638 21244 19702 21248
rect 19638 21188 19642 21244
rect 19642 21188 19698 21244
rect 19698 21188 19702 21244
rect 19638 21184 19702 21188
rect 19718 21244 19782 21248
rect 19718 21188 19722 21244
rect 19722 21188 19778 21244
rect 19778 21188 19782 21244
rect 19718 21184 19782 21188
rect 19798 21244 19862 21248
rect 19798 21188 19802 21244
rect 19802 21188 19858 21244
rect 19858 21188 19862 21244
rect 19798 21184 19862 21188
rect 50278 21244 50342 21248
rect 50278 21188 50282 21244
rect 50282 21188 50338 21244
rect 50338 21188 50342 21244
rect 50278 21184 50342 21188
rect 50358 21244 50422 21248
rect 50358 21188 50362 21244
rect 50362 21188 50418 21244
rect 50418 21188 50422 21244
rect 50358 21184 50422 21188
rect 50438 21244 50502 21248
rect 50438 21188 50442 21244
rect 50442 21188 50498 21244
rect 50498 21188 50502 21244
rect 50438 21184 50502 21188
rect 50518 21244 50582 21248
rect 50518 21188 50522 21244
rect 50522 21188 50578 21244
rect 50578 21188 50582 21244
rect 50518 21184 50582 21188
rect 4198 20700 4262 20704
rect 4198 20644 4202 20700
rect 4202 20644 4258 20700
rect 4258 20644 4262 20700
rect 4198 20640 4262 20644
rect 4278 20700 4342 20704
rect 4278 20644 4282 20700
rect 4282 20644 4338 20700
rect 4338 20644 4342 20700
rect 4278 20640 4342 20644
rect 4358 20700 4422 20704
rect 4358 20644 4362 20700
rect 4362 20644 4418 20700
rect 4418 20644 4422 20700
rect 4358 20640 4422 20644
rect 4438 20700 4502 20704
rect 4438 20644 4442 20700
rect 4442 20644 4498 20700
rect 4498 20644 4502 20700
rect 4438 20640 4502 20644
rect 34918 20700 34982 20704
rect 34918 20644 34922 20700
rect 34922 20644 34978 20700
rect 34978 20644 34982 20700
rect 34918 20640 34982 20644
rect 34998 20700 35062 20704
rect 34998 20644 35002 20700
rect 35002 20644 35058 20700
rect 35058 20644 35062 20700
rect 34998 20640 35062 20644
rect 35078 20700 35142 20704
rect 35078 20644 35082 20700
rect 35082 20644 35138 20700
rect 35138 20644 35142 20700
rect 35078 20640 35142 20644
rect 35158 20700 35222 20704
rect 35158 20644 35162 20700
rect 35162 20644 35218 20700
rect 35218 20644 35222 20700
rect 35158 20640 35222 20644
rect 19558 20156 19622 20160
rect 19558 20100 19562 20156
rect 19562 20100 19618 20156
rect 19618 20100 19622 20156
rect 19558 20096 19622 20100
rect 19638 20156 19702 20160
rect 19638 20100 19642 20156
rect 19642 20100 19698 20156
rect 19698 20100 19702 20156
rect 19638 20096 19702 20100
rect 19718 20156 19782 20160
rect 19718 20100 19722 20156
rect 19722 20100 19778 20156
rect 19778 20100 19782 20156
rect 19718 20096 19782 20100
rect 19798 20156 19862 20160
rect 19798 20100 19802 20156
rect 19802 20100 19858 20156
rect 19858 20100 19862 20156
rect 19798 20096 19862 20100
rect 50278 20156 50342 20160
rect 50278 20100 50282 20156
rect 50282 20100 50338 20156
rect 50338 20100 50342 20156
rect 50278 20096 50342 20100
rect 50358 20156 50422 20160
rect 50358 20100 50362 20156
rect 50362 20100 50418 20156
rect 50418 20100 50422 20156
rect 50358 20096 50422 20100
rect 50438 20156 50502 20160
rect 50438 20100 50442 20156
rect 50442 20100 50498 20156
rect 50498 20100 50502 20156
rect 50438 20096 50502 20100
rect 50518 20156 50582 20160
rect 50518 20100 50522 20156
rect 50522 20100 50578 20156
rect 50578 20100 50582 20156
rect 50518 20096 50582 20100
rect 4198 19612 4262 19616
rect 4198 19556 4202 19612
rect 4202 19556 4258 19612
rect 4258 19556 4262 19612
rect 4198 19552 4262 19556
rect 4278 19612 4342 19616
rect 4278 19556 4282 19612
rect 4282 19556 4338 19612
rect 4338 19556 4342 19612
rect 4278 19552 4342 19556
rect 4358 19612 4422 19616
rect 4358 19556 4362 19612
rect 4362 19556 4418 19612
rect 4418 19556 4422 19612
rect 4358 19552 4422 19556
rect 4438 19612 4502 19616
rect 4438 19556 4442 19612
rect 4442 19556 4498 19612
rect 4498 19556 4502 19612
rect 4438 19552 4502 19556
rect 34918 19612 34982 19616
rect 34918 19556 34922 19612
rect 34922 19556 34978 19612
rect 34978 19556 34982 19612
rect 34918 19552 34982 19556
rect 34998 19612 35062 19616
rect 34998 19556 35002 19612
rect 35002 19556 35058 19612
rect 35058 19556 35062 19612
rect 34998 19552 35062 19556
rect 35078 19612 35142 19616
rect 35078 19556 35082 19612
rect 35082 19556 35138 19612
rect 35138 19556 35142 19612
rect 35078 19552 35142 19556
rect 35158 19612 35222 19616
rect 35158 19556 35162 19612
rect 35162 19556 35218 19612
rect 35218 19556 35222 19612
rect 35158 19552 35222 19556
rect 19558 19068 19622 19072
rect 19558 19012 19562 19068
rect 19562 19012 19618 19068
rect 19618 19012 19622 19068
rect 19558 19008 19622 19012
rect 19638 19068 19702 19072
rect 19638 19012 19642 19068
rect 19642 19012 19698 19068
rect 19698 19012 19702 19068
rect 19638 19008 19702 19012
rect 19718 19068 19782 19072
rect 19718 19012 19722 19068
rect 19722 19012 19778 19068
rect 19778 19012 19782 19068
rect 19718 19008 19782 19012
rect 19798 19068 19862 19072
rect 19798 19012 19802 19068
rect 19802 19012 19858 19068
rect 19858 19012 19862 19068
rect 19798 19008 19862 19012
rect 50278 19068 50342 19072
rect 50278 19012 50282 19068
rect 50282 19012 50338 19068
rect 50338 19012 50342 19068
rect 50278 19008 50342 19012
rect 50358 19068 50422 19072
rect 50358 19012 50362 19068
rect 50362 19012 50418 19068
rect 50418 19012 50422 19068
rect 50358 19008 50422 19012
rect 50438 19068 50502 19072
rect 50438 19012 50442 19068
rect 50442 19012 50498 19068
rect 50498 19012 50502 19068
rect 50438 19008 50502 19012
rect 50518 19068 50582 19072
rect 50518 19012 50522 19068
rect 50522 19012 50578 19068
rect 50578 19012 50582 19068
rect 50518 19008 50582 19012
rect 4198 18524 4262 18528
rect 4198 18468 4202 18524
rect 4202 18468 4258 18524
rect 4258 18468 4262 18524
rect 4198 18464 4262 18468
rect 4278 18524 4342 18528
rect 4278 18468 4282 18524
rect 4282 18468 4338 18524
rect 4338 18468 4342 18524
rect 4278 18464 4342 18468
rect 4358 18524 4422 18528
rect 4358 18468 4362 18524
rect 4362 18468 4418 18524
rect 4418 18468 4422 18524
rect 4358 18464 4422 18468
rect 4438 18524 4502 18528
rect 4438 18468 4442 18524
rect 4442 18468 4498 18524
rect 4498 18468 4502 18524
rect 4438 18464 4502 18468
rect 34918 18524 34982 18528
rect 34918 18468 34922 18524
rect 34922 18468 34978 18524
rect 34978 18468 34982 18524
rect 34918 18464 34982 18468
rect 34998 18524 35062 18528
rect 34998 18468 35002 18524
rect 35002 18468 35058 18524
rect 35058 18468 35062 18524
rect 34998 18464 35062 18468
rect 35078 18524 35142 18528
rect 35078 18468 35082 18524
rect 35082 18468 35138 18524
rect 35138 18468 35142 18524
rect 35078 18464 35142 18468
rect 35158 18524 35222 18528
rect 35158 18468 35162 18524
rect 35162 18468 35218 18524
rect 35218 18468 35222 18524
rect 35158 18464 35222 18468
rect 19558 17980 19622 17984
rect 19558 17924 19562 17980
rect 19562 17924 19618 17980
rect 19618 17924 19622 17980
rect 19558 17920 19622 17924
rect 19638 17980 19702 17984
rect 19638 17924 19642 17980
rect 19642 17924 19698 17980
rect 19698 17924 19702 17980
rect 19638 17920 19702 17924
rect 19718 17980 19782 17984
rect 19718 17924 19722 17980
rect 19722 17924 19778 17980
rect 19778 17924 19782 17980
rect 19718 17920 19782 17924
rect 19798 17980 19862 17984
rect 19798 17924 19802 17980
rect 19802 17924 19858 17980
rect 19858 17924 19862 17980
rect 19798 17920 19862 17924
rect 50278 17980 50342 17984
rect 50278 17924 50282 17980
rect 50282 17924 50338 17980
rect 50338 17924 50342 17980
rect 50278 17920 50342 17924
rect 50358 17980 50422 17984
rect 50358 17924 50362 17980
rect 50362 17924 50418 17980
rect 50418 17924 50422 17980
rect 50358 17920 50422 17924
rect 50438 17980 50502 17984
rect 50438 17924 50442 17980
rect 50442 17924 50498 17980
rect 50498 17924 50502 17980
rect 50438 17920 50502 17924
rect 50518 17980 50582 17984
rect 50518 17924 50522 17980
rect 50522 17924 50578 17980
rect 50578 17924 50582 17980
rect 50518 17920 50582 17924
rect 4198 17436 4262 17440
rect 4198 17380 4202 17436
rect 4202 17380 4258 17436
rect 4258 17380 4262 17436
rect 4198 17376 4262 17380
rect 4278 17436 4342 17440
rect 4278 17380 4282 17436
rect 4282 17380 4338 17436
rect 4338 17380 4342 17436
rect 4278 17376 4342 17380
rect 4358 17436 4422 17440
rect 4358 17380 4362 17436
rect 4362 17380 4418 17436
rect 4418 17380 4422 17436
rect 4358 17376 4422 17380
rect 4438 17436 4502 17440
rect 4438 17380 4442 17436
rect 4442 17380 4498 17436
rect 4498 17380 4502 17436
rect 4438 17376 4502 17380
rect 34918 17436 34982 17440
rect 34918 17380 34922 17436
rect 34922 17380 34978 17436
rect 34978 17380 34982 17436
rect 34918 17376 34982 17380
rect 34998 17436 35062 17440
rect 34998 17380 35002 17436
rect 35002 17380 35058 17436
rect 35058 17380 35062 17436
rect 34998 17376 35062 17380
rect 35078 17436 35142 17440
rect 35078 17380 35082 17436
rect 35082 17380 35138 17436
rect 35138 17380 35142 17436
rect 35078 17376 35142 17380
rect 35158 17436 35222 17440
rect 35158 17380 35162 17436
rect 35162 17380 35218 17436
rect 35218 17380 35222 17436
rect 35158 17376 35222 17380
rect 19558 16892 19622 16896
rect 19558 16836 19562 16892
rect 19562 16836 19618 16892
rect 19618 16836 19622 16892
rect 19558 16832 19622 16836
rect 19638 16892 19702 16896
rect 19638 16836 19642 16892
rect 19642 16836 19698 16892
rect 19698 16836 19702 16892
rect 19638 16832 19702 16836
rect 19718 16892 19782 16896
rect 19718 16836 19722 16892
rect 19722 16836 19778 16892
rect 19778 16836 19782 16892
rect 19718 16832 19782 16836
rect 19798 16892 19862 16896
rect 19798 16836 19802 16892
rect 19802 16836 19858 16892
rect 19858 16836 19862 16892
rect 19798 16832 19862 16836
rect 50278 16892 50342 16896
rect 50278 16836 50282 16892
rect 50282 16836 50338 16892
rect 50338 16836 50342 16892
rect 50278 16832 50342 16836
rect 50358 16892 50422 16896
rect 50358 16836 50362 16892
rect 50362 16836 50418 16892
rect 50418 16836 50422 16892
rect 50358 16832 50422 16836
rect 50438 16892 50502 16896
rect 50438 16836 50442 16892
rect 50442 16836 50498 16892
rect 50498 16836 50502 16892
rect 50438 16832 50502 16836
rect 50518 16892 50582 16896
rect 50518 16836 50522 16892
rect 50522 16836 50578 16892
rect 50578 16836 50582 16892
rect 50518 16832 50582 16836
rect 4198 16348 4262 16352
rect 4198 16292 4202 16348
rect 4202 16292 4258 16348
rect 4258 16292 4262 16348
rect 4198 16288 4262 16292
rect 4278 16348 4342 16352
rect 4278 16292 4282 16348
rect 4282 16292 4338 16348
rect 4338 16292 4342 16348
rect 4278 16288 4342 16292
rect 4358 16348 4422 16352
rect 4358 16292 4362 16348
rect 4362 16292 4418 16348
rect 4418 16292 4422 16348
rect 4358 16288 4422 16292
rect 4438 16348 4502 16352
rect 4438 16292 4442 16348
rect 4442 16292 4498 16348
rect 4498 16292 4502 16348
rect 4438 16288 4502 16292
rect 34918 16348 34982 16352
rect 34918 16292 34922 16348
rect 34922 16292 34978 16348
rect 34978 16292 34982 16348
rect 34918 16288 34982 16292
rect 34998 16348 35062 16352
rect 34998 16292 35002 16348
rect 35002 16292 35058 16348
rect 35058 16292 35062 16348
rect 34998 16288 35062 16292
rect 35078 16348 35142 16352
rect 35078 16292 35082 16348
rect 35082 16292 35138 16348
rect 35138 16292 35142 16348
rect 35078 16288 35142 16292
rect 35158 16348 35222 16352
rect 35158 16292 35162 16348
rect 35162 16292 35218 16348
rect 35218 16292 35222 16348
rect 35158 16288 35222 16292
rect 19558 15804 19622 15808
rect 19558 15748 19562 15804
rect 19562 15748 19618 15804
rect 19618 15748 19622 15804
rect 19558 15744 19622 15748
rect 19638 15804 19702 15808
rect 19638 15748 19642 15804
rect 19642 15748 19698 15804
rect 19698 15748 19702 15804
rect 19638 15744 19702 15748
rect 19718 15804 19782 15808
rect 19718 15748 19722 15804
rect 19722 15748 19778 15804
rect 19778 15748 19782 15804
rect 19718 15744 19782 15748
rect 19798 15804 19862 15808
rect 19798 15748 19802 15804
rect 19802 15748 19858 15804
rect 19858 15748 19862 15804
rect 19798 15744 19862 15748
rect 50278 15804 50342 15808
rect 50278 15748 50282 15804
rect 50282 15748 50338 15804
rect 50338 15748 50342 15804
rect 50278 15744 50342 15748
rect 50358 15804 50422 15808
rect 50358 15748 50362 15804
rect 50362 15748 50418 15804
rect 50418 15748 50422 15804
rect 50358 15744 50422 15748
rect 50438 15804 50502 15808
rect 50438 15748 50442 15804
rect 50442 15748 50498 15804
rect 50498 15748 50502 15804
rect 50438 15744 50502 15748
rect 50518 15804 50582 15808
rect 50518 15748 50522 15804
rect 50522 15748 50578 15804
rect 50578 15748 50582 15804
rect 50518 15744 50582 15748
rect 4198 15260 4262 15264
rect 4198 15204 4202 15260
rect 4202 15204 4258 15260
rect 4258 15204 4262 15260
rect 4198 15200 4262 15204
rect 4278 15260 4342 15264
rect 4278 15204 4282 15260
rect 4282 15204 4338 15260
rect 4338 15204 4342 15260
rect 4278 15200 4342 15204
rect 4358 15260 4422 15264
rect 4358 15204 4362 15260
rect 4362 15204 4418 15260
rect 4418 15204 4422 15260
rect 4358 15200 4422 15204
rect 4438 15260 4502 15264
rect 4438 15204 4442 15260
rect 4442 15204 4498 15260
rect 4498 15204 4502 15260
rect 4438 15200 4502 15204
rect 34918 15260 34982 15264
rect 34918 15204 34922 15260
rect 34922 15204 34978 15260
rect 34978 15204 34982 15260
rect 34918 15200 34982 15204
rect 34998 15260 35062 15264
rect 34998 15204 35002 15260
rect 35002 15204 35058 15260
rect 35058 15204 35062 15260
rect 34998 15200 35062 15204
rect 35078 15260 35142 15264
rect 35078 15204 35082 15260
rect 35082 15204 35138 15260
rect 35138 15204 35142 15260
rect 35078 15200 35142 15204
rect 35158 15260 35222 15264
rect 35158 15204 35162 15260
rect 35162 15204 35218 15260
rect 35218 15204 35222 15260
rect 35158 15200 35222 15204
rect 23410 15132 23474 15196
rect 19558 14716 19622 14720
rect 19558 14660 19562 14716
rect 19562 14660 19618 14716
rect 19618 14660 19622 14716
rect 19558 14656 19622 14660
rect 19638 14716 19702 14720
rect 19638 14660 19642 14716
rect 19642 14660 19698 14716
rect 19698 14660 19702 14716
rect 19638 14656 19702 14660
rect 19718 14716 19782 14720
rect 19718 14660 19722 14716
rect 19722 14660 19778 14716
rect 19778 14660 19782 14716
rect 19718 14656 19782 14660
rect 19798 14716 19862 14720
rect 19798 14660 19802 14716
rect 19802 14660 19858 14716
rect 19858 14660 19862 14716
rect 19798 14656 19862 14660
rect 50278 14716 50342 14720
rect 50278 14660 50282 14716
rect 50282 14660 50338 14716
rect 50338 14660 50342 14716
rect 50278 14656 50342 14660
rect 50358 14716 50422 14720
rect 50358 14660 50362 14716
rect 50362 14660 50418 14716
rect 50418 14660 50422 14716
rect 50358 14656 50422 14660
rect 50438 14716 50502 14720
rect 50438 14660 50442 14716
rect 50442 14660 50498 14716
rect 50498 14660 50502 14716
rect 50438 14656 50502 14660
rect 50518 14716 50582 14720
rect 50518 14660 50522 14716
rect 50522 14660 50578 14716
rect 50578 14660 50582 14716
rect 50518 14656 50582 14660
rect 4198 14172 4262 14176
rect 4198 14116 4202 14172
rect 4202 14116 4258 14172
rect 4258 14116 4262 14172
rect 4198 14112 4262 14116
rect 4278 14172 4342 14176
rect 4278 14116 4282 14172
rect 4282 14116 4338 14172
rect 4338 14116 4342 14172
rect 4278 14112 4342 14116
rect 4358 14172 4422 14176
rect 4358 14116 4362 14172
rect 4362 14116 4418 14172
rect 4418 14116 4422 14172
rect 4358 14112 4422 14116
rect 4438 14172 4502 14176
rect 4438 14116 4442 14172
rect 4442 14116 4498 14172
rect 4498 14116 4502 14172
rect 4438 14112 4502 14116
rect 34918 14172 34982 14176
rect 34918 14116 34922 14172
rect 34922 14116 34978 14172
rect 34978 14116 34982 14172
rect 34918 14112 34982 14116
rect 34998 14172 35062 14176
rect 34998 14116 35002 14172
rect 35002 14116 35058 14172
rect 35058 14116 35062 14172
rect 34998 14112 35062 14116
rect 35078 14172 35142 14176
rect 35078 14116 35082 14172
rect 35082 14116 35138 14172
rect 35138 14116 35142 14172
rect 35078 14112 35142 14116
rect 35158 14172 35222 14176
rect 35158 14116 35162 14172
rect 35162 14116 35218 14172
rect 35218 14116 35222 14172
rect 35158 14112 35222 14116
rect 19558 13628 19622 13632
rect 19558 13572 19562 13628
rect 19562 13572 19618 13628
rect 19618 13572 19622 13628
rect 19558 13568 19622 13572
rect 19638 13628 19702 13632
rect 19638 13572 19642 13628
rect 19642 13572 19698 13628
rect 19698 13572 19702 13628
rect 19638 13568 19702 13572
rect 19718 13628 19782 13632
rect 19718 13572 19722 13628
rect 19722 13572 19778 13628
rect 19778 13572 19782 13628
rect 19718 13568 19782 13572
rect 19798 13628 19862 13632
rect 19798 13572 19802 13628
rect 19802 13572 19858 13628
rect 19858 13572 19862 13628
rect 19798 13568 19862 13572
rect 50278 13628 50342 13632
rect 50278 13572 50282 13628
rect 50282 13572 50338 13628
rect 50338 13572 50342 13628
rect 50278 13568 50342 13572
rect 50358 13628 50422 13632
rect 50358 13572 50362 13628
rect 50362 13572 50418 13628
rect 50418 13572 50422 13628
rect 50358 13568 50422 13572
rect 50438 13628 50502 13632
rect 50438 13572 50442 13628
rect 50442 13572 50498 13628
rect 50498 13572 50502 13628
rect 50438 13568 50502 13572
rect 50518 13628 50582 13632
rect 50518 13572 50522 13628
rect 50522 13572 50578 13628
rect 50578 13572 50582 13628
rect 50518 13568 50582 13572
rect 4198 13084 4262 13088
rect 4198 13028 4202 13084
rect 4202 13028 4258 13084
rect 4258 13028 4262 13084
rect 4198 13024 4262 13028
rect 4278 13084 4342 13088
rect 4278 13028 4282 13084
rect 4282 13028 4338 13084
rect 4338 13028 4342 13084
rect 4278 13024 4342 13028
rect 4358 13084 4422 13088
rect 4358 13028 4362 13084
rect 4362 13028 4418 13084
rect 4418 13028 4422 13084
rect 4358 13024 4422 13028
rect 4438 13084 4502 13088
rect 4438 13028 4442 13084
rect 4442 13028 4498 13084
rect 4498 13028 4502 13084
rect 4438 13024 4502 13028
rect 34918 13084 34982 13088
rect 34918 13028 34922 13084
rect 34922 13028 34978 13084
rect 34978 13028 34982 13084
rect 34918 13024 34982 13028
rect 34998 13084 35062 13088
rect 34998 13028 35002 13084
rect 35002 13028 35058 13084
rect 35058 13028 35062 13084
rect 34998 13024 35062 13028
rect 35078 13084 35142 13088
rect 35078 13028 35082 13084
rect 35082 13028 35138 13084
rect 35138 13028 35142 13084
rect 35078 13024 35142 13028
rect 35158 13084 35222 13088
rect 35158 13028 35162 13084
rect 35162 13028 35218 13084
rect 35218 13028 35222 13084
rect 35158 13024 35222 13028
rect 19558 12540 19622 12544
rect 19558 12484 19562 12540
rect 19562 12484 19618 12540
rect 19618 12484 19622 12540
rect 19558 12480 19622 12484
rect 19638 12540 19702 12544
rect 19638 12484 19642 12540
rect 19642 12484 19698 12540
rect 19698 12484 19702 12540
rect 19638 12480 19702 12484
rect 19718 12540 19782 12544
rect 19718 12484 19722 12540
rect 19722 12484 19778 12540
rect 19778 12484 19782 12540
rect 19718 12480 19782 12484
rect 19798 12540 19862 12544
rect 19798 12484 19802 12540
rect 19802 12484 19858 12540
rect 19858 12484 19862 12540
rect 19798 12480 19862 12484
rect 50278 12540 50342 12544
rect 50278 12484 50282 12540
rect 50282 12484 50338 12540
rect 50338 12484 50342 12540
rect 50278 12480 50342 12484
rect 50358 12540 50422 12544
rect 50358 12484 50362 12540
rect 50362 12484 50418 12540
rect 50418 12484 50422 12540
rect 50358 12480 50422 12484
rect 50438 12540 50502 12544
rect 50438 12484 50442 12540
rect 50442 12484 50498 12540
rect 50498 12484 50502 12540
rect 50438 12480 50502 12484
rect 50518 12540 50582 12544
rect 50518 12484 50522 12540
rect 50522 12484 50578 12540
rect 50578 12484 50582 12540
rect 50518 12480 50582 12484
rect 4198 11996 4262 12000
rect 4198 11940 4202 11996
rect 4202 11940 4258 11996
rect 4258 11940 4262 11996
rect 4198 11936 4262 11940
rect 4278 11996 4342 12000
rect 4278 11940 4282 11996
rect 4282 11940 4338 11996
rect 4338 11940 4342 11996
rect 4278 11936 4342 11940
rect 4358 11996 4422 12000
rect 4358 11940 4362 11996
rect 4362 11940 4418 11996
rect 4418 11940 4422 11996
rect 4358 11936 4422 11940
rect 4438 11996 4502 12000
rect 4438 11940 4442 11996
rect 4442 11940 4498 11996
rect 4498 11940 4502 11996
rect 4438 11936 4502 11940
rect 34918 11996 34982 12000
rect 34918 11940 34922 11996
rect 34922 11940 34978 11996
rect 34978 11940 34982 11996
rect 34918 11936 34982 11940
rect 34998 11996 35062 12000
rect 34998 11940 35002 11996
rect 35002 11940 35058 11996
rect 35058 11940 35062 11996
rect 34998 11936 35062 11940
rect 35078 11996 35142 12000
rect 35078 11940 35082 11996
rect 35082 11940 35138 11996
rect 35138 11940 35142 11996
rect 35078 11936 35142 11940
rect 35158 11996 35222 12000
rect 35158 11940 35162 11996
rect 35162 11940 35218 11996
rect 35218 11940 35222 11996
rect 35158 11936 35222 11940
rect 19558 11452 19622 11456
rect 19558 11396 19562 11452
rect 19562 11396 19618 11452
rect 19618 11396 19622 11452
rect 19558 11392 19622 11396
rect 19638 11452 19702 11456
rect 19638 11396 19642 11452
rect 19642 11396 19698 11452
rect 19698 11396 19702 11452
rect 19638 11392 19702 11396
rect 19718 11452 19782 11456
rect 19718 11396 19722 11452
rect 19722 11396 19778 11452
rect 19778 11396 19782 11452
rect 19718 11392 19782 11396
rect 19798 11452 19862 11456
rect 19798 11396 19802 11452
rect 19802 11396 19858 11452
rect 19858 11396 19862 11452
rect 19798 11392 19862 11396
rect 50278 11452 50342 11456
rect 50278 11396 50282 11452
rect 50282 11396 50338 11452
rect 50338 11396 50342 11452
rect 50278 11392 50342 11396
rect 50358 11452 50422 11456
rect 50358 11396 50362 11452
rect 50362 11396 50418 11452
rect 50418 11396 50422 11452
rect 50358 11392 50422 11396
rect 50438 11452 50502 11456
rect 50438 11396 50442 11452
rect 50442 11396 50498 11452
rect 50498 11396 50502 11452
rect 50438 11392 50502 11396
rect 50518 11452 50582 11456
rect 50518 11396 50522 11452
rect 50522 11396 50578 11452
rect 50578 11396 50582 11452
rect 50518 11392 50582 11396
rect 4198 10908 4262 10912
rect 4198 10852 4202 10908
rect 4202 10852 4258 10908
rect 4258 10852 4262 10908
rect 4198 10848 4262 10852
rect 4278 10908 4342 10912
rect 4278 10852 4282 10908
rect 4282 10852 4338 10908
rect 4338 10852 4342 10908
rect 4278 10848 4342 10852
rect 4358 10908 4422 10912
rect 4358 10852 4362 10908
rect 4362 10852 4418 10908
rect 4418 10852 4422 10908
rect 4358 10848 4422 10852
rect 4438 10908 4502 10912
rect 4438 10852 4442 10908
rect 4442 10852 4498 10908
rect 4498 10852 4502 10908
rect 4438 10848 4502 10852
rect 34918 10908 34982 10912
rect 34918 10852 34922 10908
rect 34922 10852 34978 10908
rect 34978 10852 34982 10908
rect 34918 10848 34982 10852
rect 34998 10908 35062 10912
rect 34998 10852 35002 10908
rect 35002 10852 35058 10908
rect 35058 10852 35062 10908
rect 34998 10848 35062 10852
rect 35078 10908 35142 10912
rect 35078 10852 35082 10908
rect 35082 10852 35138 10908
rect 35138 10852 35142 10908
rect 35078 10848 35142 10852
rect 35158 10908 35222 10912
rect 35158 10852 35162 10908
rect 35162 10852 35218 10908
rect 35218 10852 35222 10908
rect 35158 10848 35222 10852
rect 19558 10364 19622 10368
rect 19558 10308 19562 10364
rect 19562 10308 19618 10364
rect 19618 10308 19622 10364
rect 19558 10304 19622 10308
rect 19638 10364 19702 10368
rect 19638 10308 19642 10364
rect 19642 10308 19698 10364
rect 19698 10308 19702 10364
rect 19638 10304 19702 10308
rect 19718 10364 19782 10368
rect 19718 10308 19722 10364
rect 19722 10308 19778 10364
rect 19778 10308 19782 10364
rect 19718 10304 19782 10308
rect 19798 10364 19862 10368
rect 19798 10308 19802 10364
rect 19802 10308 19858 10364
rect 19858 10308 19862 10364
rect 19798 10304 19862 10308
rect 50278 10364 50342 10368
rect 50278 10308 50282 10364
rect 50282 10308 50338 10364
rect 50338 10308 50342 10364
rect 50278 10304 50342 10308
rect 50358 10364 50422 10368
rect 50358 10308 50362 10364
rect 50362 10308 50418 10364
rect 50418 10308 50422 10364
rect 50358 10304 50422 10308
rect 50438 10364 50502 10368
rect 50438 10308 50442 10364
rect 50442 10308 50498 10364
rect 50498 10308 50502 10364
rect 50438 10304 50502 10308
rect 50518 10364 50582 10368
rect 50518 10308 50522 10364
rect 50522 10308 50578 10364
rect 50578 10308 50582 10364
rect 50518 10304 50582 10308
rect 4198 9820 4262 9824
rect 4198 9764 4202 9820
rect 4202 9764 4258 9820
rect 4258 9764 4262 9820
rect 4198 9760 4262 9764
rect 4278 9820 4342 9824
rect 4278 9764 4282 9820
rect 4282 9764 4338 9820
rect 4338 9764 4342 9820
rect 4278 9760 4342 9764
rect 4358 9820 4422 9824
rect 4358 9764 4362 9820
rect 4362 9764 4418 9820
rect 4418 9764 4422 9820
rect 4358 9760 4422 9764
rect 4438 9820 4502 9824
rect 4438 9764 4442 9820
rect 4442 9764 4498 9820
rect 4498 9764 4502 9820
rect 4438 9760 4502 9764
rect 34918 9820 34982 9824
rect 34918 9764 34922 9820
rect 34922 9764 34978 9820
rect 34978 9764 34982 9820
rect 34918 9760 34982 9764
rect 34998 9820 35062 9824
rect 34998 9764 35002 9820
rect 35002 9764 35058 9820
rect 35058 9764 35062 9820
rect 34998 9760 35062 9764
rect 35078 9820 35142 9824
rect 35078 9764 35082 9820
rect 35082 9764 35138 9820
rect 35138 9764 35142 9820
rect 35078 9760 35142 9764
rect 35158 9820 35222 9824
rect 35158 9764 35162 9820
rect 35162 9764 35218 9820
rect 35218 9764 35222 9820
rect 35158 9760 35222 9764
rect 19558 9276 19622 9280
rect 19558 9220 19562 9276
rect 19562 9220 19618 9276
rect 19618 9220 19622 9276
rect 19558 9216 19622 9220
rect 19638 9276 19702 9280
rect 19638 9220 19642 9276
rect 19642 9220 19698 9276
rect 19698 9220 19702 9276
rect 19638 9216 19702 9220
rect 19718 9276 19782 9280
rect 19718 9220 19722 9276
rect 19722 9220 19778 9276
rect 19778 9220 19782 9276
rect 19718 9216 19782 9220
rect 19798 9276 19862 9280
rect 19798 9220 19802 9276
rect 19802 9220 19858 9276
rect 19858 9220 19862 9276
rect 19798 9216 19862 9220
rect 50278 9276 50342 9280
rect 50278 9220 50282 9276
rect 50282 9220 50338 9276
rect 50338 9220 50342 9276
rect 50278 9216 50342 9220
rect 50358 9276 50422 9280
rect 50358 9220 50362 9276
rect 50362 9220 50418 9276
rect 50418 9220 50422 9276
rect 50358 9216 50422 9220
rect 50438 9276 50502 9280
rect 50438 9220 50442 9276
rect 50442 9220 50498 9276
rect 50498 9220 50502 9276
rect 50438 9216 50502 9220
rect 50518 9276 50582 9280
rect 50518 9220 50522 9276
rect 50522 9220 50578 9276
rect 50578 9220 50582 9276
rect 50518 9216 50582 9220
rect 4198 8732 4262 8736
rect 4198 8676 4202 8732
rect 4202 8676 4258 8732
rect 4258 8676 4262 8732
rect 4198 8672 4262 8676
rect 4278 8732 4342 8736
rect 4278 8676 4282 8732
rect 4282 8676 4338 8732
rect 4338 8676 4342 8732
rect 4278 8672 4342 8676
rect 4358 8732 4422 8736
rect 4358 8676 4362 8732
rect 4362 8676 4418 8732
rect 4418 8676 4422 8732
rect 4358 8672 4422 8676
rect 4438 8732 4502 8736
rect 4438 8676 4442 8732
rect 4442 8676 4498 8732
rect 4498 8676 4502 8732
rect 4438 8672 4502 8676
rect 34918 8732 34982 8736
rect 34918 8676 34922 8732
rect 34922 8676 34978 8732
rect 34978 8676 34982 8732
rect 34918 8672 34982 8676
rect 34998 8732 35062 8736
rect 34998 8676 35002 8732
rect 35002 8676 35058 8732
rect 35058 8676 35062 8732
rect 34998 8672 35062 8676
rect 35078 8732 35142 8736
rect 35078 8676 35082 8732
rect 35082 8676 35138 8732
rect 35138 8676 35142 8732
rect 35078 8672 35142 8676
rect 35158 8732 35222 8736
rect 35158 8676 35162 8732
rect 35162 8676 35218 8732
rect 35218 8676 35222 8732
rect 35158 8672 35222 8676
rect 19558 8188 19622 8192
rect 19558 8132 19562 8188
rect 19562 8132 19618 8188
rect 19618 8132 19622 8188
rect 19558 8128 19622 8132
rect 19638 8188 19702 8192
rect 19638 8132 19642 8188
rect 19642 8132 19698 8188
rect 19698 8132 19702 8188
rect 19638 8128 19702 8132
rect 19718 8188 19782 8192
rect 19718 8132 19722 8188
rect 19722 8132 19778 8188
rect 19778 8132 19782 8188
rect 19718 8128 19782 8132
rect 19798 8188 19862 8192
rect 19798 8132 19802 8188
rect 19802 8132 19858 8188
rect 19858 8132 19862 8188
rect 19798 8128 19862 8132
rect 50278 8188 50342 8192
rect 50278 8132 50282 8188
rect 50282 8132 50338 8188
rect 50338 8132 50342 8188
rect 50278 8128 50342 8132
rect 50358 8188 50422 8192
rect 50358 8132 50362 8188
rect 50362 8132 50418 8188
rect 50418 8132 50422 8188
rect 50358 8128 50422 8132
rect 50438 8188 50502 8192
rect 50438 8132 50442 8188
rect 50442 8132 50498 8188
rect 50498 8132 50502 8188
rect 50438 8128 50502 8132
rect 50518 8188 50582 8192
rect 50518 8132 50522 8188
rect 50522 8132 50578 8188
rect 50578 8132 50582 8188
rect 50518 8128 50582 8132
rect 20282 7652 20346 7716
rect 4198 7644 4262 7648
rect 4198 7588 4202 7644
rect 4202 7588 4258 7644
rect 4258 7588 4262 7644
rect 4198 7584 4262 7588
rect 4278 7644 4342 7648
rect 4278 7588 4282 7644
rect 4282 7588 4338 7644
rect 4338 7588 4342 7644
rect 4278 7584 4342 7588
rect 4358 7644 4422 7648
rect 4358 7588 4362 7644
rect 4362 7588 4418 7644
rect 4418 7588 4422 7644
rect 4358 7584 4422 7588
rect 4438 7644 4502 7648
rect 4438 7588 4442 7644
rect 4442 7588 4498 7644
rect 4498 7588 4502 7644
rect 4438 7584 4502 7588
rect 34918 7644 34982 7648
rect 34918 7588 34922 7644
rect 34922 7588 34978 7644
rect 34978 7588 34982 7644
rect 34918 7584 34982 7588
rect 34998 7644 35062 7648
rect 34998 7588 35002 7644
rect 35002 7588 35058 7644
rect 35058 7588 35062 7644
rect 34998 7584 35062 7588
rect 35078 7644 35142 7648
rect 35078 7588 35082 7644
rect 35082 7588 35138 7644
rect 35138 7588 35142 7644
rect 35078 7584 35142 7588
rect 35158 7644 35222 7648
rect 35158 7588 35162 7644
rect 35162 7588 35218 7644
rect 35218 7588 35222 7644
rect 35158 7584 35222 7588
rect 19558 7100 19622 7104
rect 19558 7044 19562 7100
rect 19562 7044 19618 7100
rect 19618 7044 19622 7100
rect 19558 7040 19622 7044
rect 19638 7100 19702 7104
rect 19638 7044 19642 7100
rect 19642 7044 19698 7100
rect 19698 7044 19702 7100
rect 19638 7040 19702 7044
rect 19718 7100 19782 7104
rect 19718 7044 19722 7100
rect 19722 7044 19778 7100
rect 19778 7044 19782 7100
rect 19718 7040 19782 7044
rect 19798 7100 19862 7104
rect 19798 7044 19802 7100
rect 19802 7044 19858 7100
rect 19858 7044 19862 7100
rect 19798 7040 19862 7044
rect 50278 7100 50342 7104
rect 50278 7044 50282 7100
rect 50282 7044 50338 7100
rect 50338 7044 50342 7100
rect 50278 7040 50342 7044
rect 50358 7100 50422 7104
rect 50358 7044 50362 7100
rect 50362 7044 50418 7100
rect 50418 7044 50422 7100
rect 50358 7040 50422 7044
rect 50438 7100 50502 7104
rect 50438 7044 50442 7100
rect 50442 7044 50498 7100
rect 50498 7044 50502 7100
rect 50438 7040 50502 7044
rect 50518 7100 50582 7104
rect 50518 7044 50522 7100
rect 50522 7044 50578 7100
rect 50578 7044 50582 7100
rect 50518 7040 50582 7044
rect 4198 6556 4262 6560
rect 4198 6500 4202 6556
rect 4202 6500 4258 6556
rect 4258 6500 4262 6556
rect 4198 6496 4262 6500
rect 4278 6556 4342 6560
rect 4278 6500 4282 6556
rect 4282 6500 4338 6556
rect 4338 6500 4342 6556
rect 4278 6496 4342 6500
rect 4358 6556 4422 6560
rect 4358 6500 4362 6556
rect 4362 6500 4418 6556
rect 4418 6500 4422 6556
rect 4358 6496 4422 6500
rect 4438 6556 4502 6560
rect 4438 6500 4442 6556
rect 4442 6500 4498 6556
rect 4498 6500 4502 6556
rect 4438 6496 4502 6500
rect 34918 6556 34982 6560
rect 34918 6500 34922 6556
rect 34922 6500 34978 6556
rect 34978 6500 34982 6556
rect 34918 6496 34982 6500
rect 34998 6556 35062 6560
rect 34998 6500 35002 6556
rect 35002 6500 35058 6556
rect 35058 6500 35062 6556
rect 34998 6496 35062 6500
rect 35078 6556 35142 6560
rect 35078 6500 35082 6556
rect 35082 6500 35138 6556
rect 35138 6500 35142 6556
rect 35078 6496 35142 6500
rect 35158 6556 35222 6560
rect 35158 6500 35162 6556
rect 35162 6500 35218 6556
rect 35218 6500 35222 6556
rect 35158 6496 35222 6500
rect 19558 6012 19622 6016
rect 19558 5956 19562 6012
rect 19562 5956 19618 6012
rect 19618 5956 19622 6012
rect 19558 5952 19622 5956
rect 19638 6012 19702 6016
rect 19638 5956 19642 6012
rect 19642 5956 19698 6012
rect 19698 5956 19702 6012
rect 19638 5952 19702 5956
rect 19718 6012 19782 6016
rect 19718 5956 19722 6012
rect 19722 5956 19778 6012
rect 19778 5956 19782 6012
rect 19718 5952 19782 5956
rect 19798 6012 19862 6016
rect 19798 5956 19802 6012
rect 19802 5956 19858 6012
rect 19858 5956 19862 6012
rect 19798 5952 19862 5956
rect 50278 6012 50342 6016
rect 50278 5956 50282 6012
rect 50282 5956 50338 6012
rect 50338 5956 50342 6012
rect 50278 5952 50342 5956
rect 50358 6012 50422 6016
rect 50358 5956 50362 6012
rect 50362 5956 50418 6012
rect 50418 5956 50422 6012
rect 50358 5952 50422 5956
rect 50438 6012 50502 6016
rect 50438 5956 50442 6012
rect 50442 5956 50498 6012
rect 50498 5956 50502 6012
rect 50438 5952 50502 5956
rect 50518 6012 50582 6016
rect 50518 5956 50522 6012
rect 50522 5956 50578 6012
rect 50578 5956 50582 6012
rect 50518 5952 50582 5956
rect 4198 5468 4262 5472
rect 4198 5412 4202 5468
rect 4202 5412 4258 5468
rect 4258 5412 4262 5468
rect 4198 5408 4262 5412
rect 4278 5468 4342 5472
rect 4278 5412 4282 5468
rect 4282 5412 4338 5468
rect 4338 5412 4342 5468
rect 4278 5408 4342 5412
rect 4358 5468 4422 5472
rect 4358 5412 4362 5468
rect 4362 5412 4418 5468
rect 4418 5412 4422 5468
rect 4358 5408 4422 5412
rect 4438 5468 4502 5472
rect 4438 5412 4442 5468
rect 4442 5412 4498 5468
rect 4498 5412 4502 5468
rect 4438 5408 4502 5412
rect 34918 5468 34982 5472
rect 34918 5412 34922 5468
rect 34922 5412 34978 5468
rect 34978 5412 34982 5468
rect 34918 5408 34982 5412
rect 34998 5468 35062 5472
rect 34998 5412 35002 5468
rect 35002 5412 35058 5468
rect 35058 5412 35062 5468
rect 34998 5408 35062 5412
rect 35078 5468 35142 5472
rect 35078 5412 35082 5468
rect 35082 5412 35138 5468
rect 35138 5412 35142 5468
rect 35078 5408 35142 5412
rect 35158 5468 35222 5472
rect 35158 5412 35162 5468
rect 35162 5412 35218 5468
rect 35218 5412 35222 5468
rect 35158 5408 35222 5412
rect 19558 4924 19622 4928
rect 19558 4868 19562 4924
rect 19562 4868 19618 4924
rect 19618 4868 19622 4924
rect 19558 4864 19622 4868
rect 19638 4924 19702 4928
rect 19638 4868 19642 4924
rect 19642 4868 19698 4924
rect 19698 4868 19702 4924
rect 19638 4864 19702 4868
rect 19718 4924 19782 4928
rect 19718 4868 19722 4924
rect 19722 4868 19778 4924
rect 19778 4868 19782 4924
rect 19718 4864 19782 4868
rect 19798 4924 19862 4928
rect 19798 4868 19802 4924
rect 19802 4868 19858 4924
rect 19858 4868 19862 4924
rect 19798 4864 19862 4868
rect 50278 4924 50342 4928
rect 50278 4868 50282 4924
rect 50282 4868 50338 4924
rect 50338 4868 50342 4924
rect 50278 4864 50342 4868
rect 50358 4924 50422 4928
rect 50358 4868 50362 4924
rect 50362 4868 50418 4924
rect 50418 4868 50422 4924
rect 50358 4864 50422 4868
rect 50438 4924 50502 4928
rect 50438 4868 50442 4924
rect 50442 4868 50498 4924
rect 50498 4868 50502 4924
rect 50438 4864 50502 4868
rect 50518 4924 50582 4928
rect 50518 4868 50522 4924
rect 50522 4868 50578 4924
rect 50578 4868 50582 4924
rect 50518 4864 50582 4868
rect 4198 4380 4262 4384
rect 4198 4324 4202 4380
rect 4202 4324 4258 4380
rect 4258 4324 4262 4380
rect 4198 4320 4262 4324
rect 4278 4380 4342 4384
rect 4278 4324 4282 4380
rect 4282 4324 4338 4380
rect 4338 4324 4342 4380
rect 4278 4320 4342 4324
rect 4358 4380 4422 4384
rect 4358 4324 4362 4380
rect 4362 4324 4418 4380
rect 4418 4324 4422 4380
rect 4358 4320 4422 4324
rect 4438 4380 4502 4384
rect 4438 4324 4442 4380
rect 4442 4324 4498 4380
rect 4498 4324 4502 4380
rect 4438 4320 4502 4324
rect 34918 4380 34982 4384
rect 34918 4324 34922 4380
rect 34922 4324 34978 4380
rect 34978 4324 34982 4380
rect 34918 4320 34982 4324
rect 34998 4380 35062 4384
rect 34998 4324 35002 4380
rect 35002 4324 35058 4380
rect 35058 4324 35062 4380
rect 34998 4320 35062 4324
rect 35078 4380 35142 4384
rect 35078 4324 35082 4380
rect 35082 4324 35138 4380
rect 35138 4324 35142 4380
rect 35078 4320 35142 4324
rect 35158 4380 35222 4384
rect 35158 4324 35162 4380
rect 35162 4324 35218 4380
rect 35218 4324 35222 4380
rect 35158 4320 35222 4324
rect 19558 3836 19622 3840
rect 19558 3780 19562 3836
rect 19562 3780 19618 3836
rect 19618 3780 19622 3836
rect 19558 3776 19622 3780
rect 19638 3836 19702 3840
rect 19638 3780 19642 3836
rect 19642 3780 19698 3836
rect 19698 3780 19702 3836
rect 19638 3776 19702 3780
rect 19718 3836 19782 3840
rect 19718 3780 19722 3836
rect 19722 3780 19778 3836
rect 19778 3780 19782 3836
rect 19718 3776 19782 3780
rect 19798 3836 19862 3840
rect 19798 3780 19802 3836
rect 19802 3780 19858 3836
rect 19858 3780 19862 3836
rect 19798 3776 19862 3780
rect 41258 3844 41322 3908
rect 50278 3836 50342 3840
rect 50278 3780 50282 3836
rect 50282 3780 50338 3836
rect 50338 3780 50342 3836
rect 50278 3776 50342 3780
rect 50358 3836 50422 3840
rect 50358 3780 50362 3836
rect 50362 3780 50418 3836
rect 50418 3780 50422 3836
rect 50358 3776 50422 3780
rect 50438 3836 50502 3840
rect 50438 3780 50442 3836
rect 50442 3780 50498 3836
rect 50498 3780 50502 3836
rect 50438 3776 50502 3780
rect 50518 3836 50582 3840
rect 50518 3780 50522 3836
rect 50522 3780 50578 3836
rect 50578 3780 50582 3836
rect 50518 3776 50582 3780
rect 4198 3292 4262 3296
rect 4198 3236 4202 3292
rect 4202 3236 4258 3292
rect 4258 3236 4262 3292
rect 4198 3232 4262 3236
rect 4278 3292 4342 3296
rect 4278 3236 4282 3292
rect 4282 3236 4338 3292
rect 4338 3236 4342 3292
rect 4278 3232 4342 3236
rect 4358 3292 4422 3296
rect 4358 3236 4362 3292
rect 4362 3236 4418 3292
rect 4418 3236 4422 3292
rect 4358 3232 4422 3236
rect 4438 3292 4502 3296
rect 4438 3236 4442 3292
rect 4442 3236 4498 3292
rect 4498 3236 4502 3292
rect 4438 3232 4502 3236
rect 34918 3292 34982 3296
rect 34918 3236 34922 3292
rect 34922 3236 34978 3292
rect 34978 3236 34982 3292
rect 34918 3232 34982 3236
rect 34998 3292 35062 3296
rect 34998 3236 35002 3292
rect 35002 3236 35058 3292
rect 35058 3236 35062 3292
rect 34998 3232 35062 3236
rect 35078 3292 35142 3296
rect 35078 3236 35082 3292
rect 35082 3236 35138 3292
rect 35138 3236 35142 3292
rect 35078 3232 35142 3236
rect 35158 3292 35222 3296
rect 35158 3236 35162 3292
rect 35162 3236 35218 3292
rect 35218 3236 35222 3292
rect 35158 3232 35222 3236
rect 41258 2892 41322 2956
rect 19558 2748 19622 2752
rect 19558 2692 19562 2748
rect 19562 2692 19618 2748
rect 19618 2692 19622 2748
rect 19558 2688 19622 2692
rect 19638 2748 19702 2752
rect 19638 2692 19642 2748
rect 19642 2692 19698 2748
rect 19698 2692 19702 2748
rect 19638 2688 19702 2692
rect 19718 2748 19782 2752
rect 19718 2692 19722 2748
rect 19722 2692 19778 2748
rect 19778 2692 19782 2748
rect 19718 2688 19782 2692
rect 19798 2748 19862 2752
rect 19798 2692 19802 2748
rect 19802 2692 19858 2748
rect 19858 2692 19862 2748
rect 19798 2688 19862 2692
rect 50278 2748 50342 2752
rect 50278 2692 50282 2748
rect 50282 2692 50338 2748
rect 50338 2692 50342 2748
rect 50278 2688 50342 2692
rect 50358 2748 50422 2752
rect 50358 2692 50362 2748
rect 50362 2692 50418 2748
rect 50418 2692 50422 2748
rect 50358 2688 50422 2692
rect 50438 2748 50502 2752
rect 50438 2692 50442 2748
rect 50442 2692 50498 2748
rect 50498 2692 50502 2748
rect 50438 2688 50502 2692
rect 50518 2748 50582 2752
rect 50518 2692 50522 2748
rect 50522 2692 50578 2748
rect 50578 2692 50582 2748
rect 50518 2688 50582 2692
rect 4198 2204 4262 2208
rect 4198 2148 4202 2204
rect 4202 2148 4258 2204
rect 4258 2148 4262 2204
rect 4198 2144 4262 2148
rect 4278 2204 4342 2208
rect 4278 2148 4282 2204
rect 4282 2148 4338 2204
rect 4338 2148 4342 2204
rect 4278 2144 4342 2148
rect 4358 2204 4422 2208
rect 4358 2148 4362 2204
rect 4362 2148 4418 2204
rect 4418 2148 4422 2204
rect 4358 2144 4422 2148
rect 4438 2204 4502 2208
rect 4438 2148 4442 2204
rect 4442 2148 4498 2204
rect 4498 2148 4502 2204
rect 4438 2144 4502 2148
rect 34918 2204 34982 2208
rect 34918 2148 34922 2204
rect 34922 2148 34978 2204
rect 34978 2148 34982 2204
rect 34918 2144 34982 2148
rect 34998 2204 35062 2208
rect 34998 2148 35002 2204
rect 35002 2148 35058 2204
rect 35058 2148 35062 2204
rect 34998 2144 35062 2148
rect 35078 2204 35142 2208
rect 35078 2148 35082 2204
rect 35082 2148 35138 2204
rect 35138 2148 35142 2204
rect 35078 2144 35142 2148
rect 35158 2204 35222 2208
rect 35158 2148 35162 2204
rect 35162 2148 35218 2204
rect 35218 2148 35222 2204
rect 35158 2144 35222 2148
rect 20282 852 20346 916
<< metal4 >>
rect 4190 57696 4510 57712
rect 4190 57632 4198 57696
rect 4262 57632 4278 57696
rect 4342 57632 4358 57696
rect 4422 57632 4438 57696
rect 4502 57632 4510 57696
rect 4190 56608 4510 57632
rect 4190 56544 4198 56608
rect 4262 56544 4278 56608
rect 4342 56544 4358 56608
rect 4422 56544 4438 56608
rect 4502 56544 4510 56608
rect 4190 55520 4510 56544
rect 4190 55456 4198 55520
rect 4262 55456 4278 55520
rect 4342 55456 4358 55520
rect 4422 55456 4438 55520
rect 4502 55456 4510 55520
rect 4190 54432 4510 55456
rect 4190 54368 4198 54432
rect 4262 54368 4278 54432
rect 4342 54368 4358 54432
rect 4422 54368 4438 54432
rect 4502 54368 4510 54432
rect 4190 53344 4510 54368
rect 4190 53280 4198 53344
rect 4262 53280 4278 53344
rect 4342 53280 4358 53344
rect 4422 53280 4438 53344
rect 4502 53280 4510 53344
rect 4190 52256 4510 53280
rect 4190 52192 4198 52256
rect 4262 52192 4278 52256
rect 4342 52192 4358 52256
rect 4422 52192 4438 52256
rect 4502 52192 4510 52256
rect 4190 51168 4510 52192
rect 4190 51104 4198 51168
rect 4262 51104 4278 51168
rect 4342 51104 4358 51168
rect 4422 51104 4438 51168
rect 4502 51104 4510 51168
rect 4190 50080 4510 51104
rect 4190 50016 4198 50080
rect 4262 50016 4278 50080
rect 4342 50016 4358 50080
rect 4422 50016 4438 50080
rect 4502 50016 4510 50080
rect 4190 48992 4510 50016
rect 4190 48928 4198 48992
rect 4262 48928 4278 48992
rect 4342 48928 4358 48992
rect 4422 48928 4438 48992
rect 4502 48928 4510 48992
rect 4190 47904 4510 48928
rect 4190 47840 4198 47904
rect 4262 47840 4278 47904
rect 4342 47840 4358 47904
rect 4422 47840 4438 47904
rect 4502 47840 4510 47904
rect 4190 46816 4510 47840
rect 4190 46752 4198 46816
rect 4262 46752 4278 46816
rect 4342 46752 4358 46816
rect 4422 46752 4438 46816
rect 4502 46752 4510 46816
rect 4190 45728 4510 46752
rect 4190 45664 4198 45728
rect 4262 45664 4278 45728
rect 4342 45664 4358 45728
rect 4422 45664 4438 45728
rect 4502 45664 4510 45728
rect 4190 44640 4510 45664
rect 4190 44576 4198 44640
rect 4262 44576 4278 44640
rect 4342 44576 4358 44640
rect 4422 44576 4438 44640
rect 4502 44576 4510 44640
rect 4190 43552 4510 44576
rect 4190 43488 4198 43552
rect 4262 43488 4278 43552
rect 4342 43488 4358 43552
rect 4422 43488 4438 43552
rect 4502 43488 4510 43552
rect 4190 42464 4510 43488
rect 4190 42400 4198 42464
rect 4262 42400 4278 42464
rect 4342 42400 4358 42464
rect 4422 42400 4438 42464
rect 4502 42400 4510 42464
rect 4190 41376 4510 42400
rect 4190 41312 4198 41376
rect 4262 41312 4278 41376
rect 4342 41312 4358 41376
rect 4422 41312 4438 41376
rect 4502 41312 4510 41376
rect 4190 40288 4510 41312
rect 4190 40224 4198 40288
rect 4262 40224 4278 40288
rect 4342 40224 4358 40288
rect 4422 40224 4438 40288
rect 4502 40224 4510 40288
rect 4190 39200 4510 40224
rect 4190 39136 4198 39200
rect 4262 39136 4278 39200
rect 4342 39136 4358 39200
rect 4422 39136 4438 39200
rect 4502 39136 4510 39200
rect 4190 38112 4510 39136
rect 4190 38048 4198 38112
rect 4262 38048 4278 38112
rect 4342 38048 4358 38112
rect 4422 38048 4438 38112
rect 4502 38048 4510 38112
rect 4190 37024 4510 38048
rect 4190 36960 4198 37024
rect 4262 36960 4278 37024
rect 4342 36960 4358 37024
rect 4422 36960 4438 37024
rect 4502 36960 4510 37024
rect 4190 35936 4510 36960
rect 4190 35872 4198 35936
rect 4262 35872 4278 35936
rect 4342 35872 4358 35936
rect 4422 35872 4438 35936
rect 4502 35872 4510 35936
rect 4190 34848 4510 35872
rect 4190 34784 4198 34848
rect 4262 34784 4278 34848
rect 4342 34784 4358 34848
rect 4422 34784 4438 34848
rect 4502 34784 4510 34848
rect 4190 33760 4510 34784
rect 4190 33696 4198 33760
rect 4262 33696 4278 33760
rect 4342 33696 4358 33760
rect 4422 33696 4438 33760
rect 4502 33696 4510 33760
rect 4190 32672 4510 33696
rect 4190 32608 4198 32672
rect 4262 32608 4278 32672
rect 4342 32608 4358 32672
rect 4422 32608 4438 32672
rect 4502 32608 4510 32672
rect 4190 31584 4510 32608
rect 4190 31520 4198 31584
rect 4262 31520 4278 31584
rect 4342 31520 4358 31584
rect 4422 31520 4438 31584
rect 4502 31520 4510 31584
rect 4190 30496 4510 31520
rect 4190 30432 4198 30496
rect 4262 30432 4278 30496
rect 4342 30432 4358 30496
rect 4422 30432 4438 30496
rect 4502 30432 4510 30496
rect 4190 29408 4510 30432
rect 4190 29344 4198 29408
rect 4262 29344 4278 29408
rect 4342 29344 4358 29408
rect 4422 29344 4438 29408
rect 4502 29344 4510 29408
rect 4190 28320 4510 29344
rect 4190 28256 4198 28320
rect 4262 28256 4278 28320
rect 4342 28256 4358 28320
rect 4422 28256 4438 28320
rect 4502 28256 4510 28320
rect 4190 27232 4510 28256
rect 4190 27168 4198 27232
rect 4262 27168 4278 27232
rect 4342 27168 4358 27232
rect 4422 27168 4438 27232
rect 4502 27168 4510 27232
rect 4190 26144 4510 27168
rect 4190 26080 4198 26144
rect 4262 26080 4278 26144
rect 4342 26080 4358 26144
rect 4422 26080 4438 26144
rect 4502 26080 4510 26144
rect 4190 25056 4510 26080
rect 4190 24992 4198 25056
rect 4262 24992 4278 25056
rect 4342 24992 4358 25056
rect 4422 24992 4438 25056
rect 4502 24992 4510 25056
rect 4190 23968 4510 24992
rect 4190 23904 4198 23968
rect 4262 23904 4278 23968
rect 4342 23904 4358 23968
rect 4422 23904 4438 23968
rect 4502 23904 4510 23968
rect 4190 22880 4510 23904
rect 4190 22816 4198 22880
rect 4262 22816 4278 22880
rect 4342 22816 4358 22880
rect 4422 22816 4438 22880
rect 4502 22816 4510 22880
rect 4190 21792 4510 22816
rect 4190 21728 4198 21792
rect 4262 21728 4278 21792
rect 4342 21728 4358 21792
rect 4422 21728 4438 21792
rect 4502 21728 4510 21792
rect 4190 20704 4510 21728
rect 4190 20640 4198 20704
rect 4262 20640 4278 20704
rect 4342 20640 4358 20704
rect 4422 20640 4438 20704
rect 4502 20640 4510 20704
rect 4190 19616 4510 20640
rect 4190 19552 4198 19616
rect 4262 19552 4278 19616
rect 4342 19552 4358 19616
rect 4422 19552 4438 19616
rect 4502 19552 4510 19616
rect 4190 18528 4510 19552
rect 4190 18464 4198 18528
rect 4262 18464 4278 18528
rect 4342 18464 4358 18528
rect 4422 18464 4438 18528
rect 4502 18464 4510 18528
rect 4190 17440 4510 18464
rect 4190 17376 4198 17440
rect 4262 17376 4278 17440
rect 4342 17376 4358 17440
rect 4422 17376 4438 17440
rect 4502 17376 4510 17440
rect 4190 16352 4510 17376
rect 4190 16288 4198 16352
rect 4262 16288 4278 16352
rect 4342 16288 4358 16352
rect 4422 16288 4438 16352
rect 4502 16288 4510 16352
rect 4190 15264 4510 16288
rect 4190 15200 4198 15264
rect 4262 15200 4278 15264
rect 4342 15200 4358 15264
rect 4422 15200 4438 15264
rect 4502 15200 4510 15264
rect 4190 14176 4510 15200
rect 4190 14112 4198 14176
rect 4262 14112 4278 14176
rect 4342 14112 4358 14176
rect 4422 14112 4438 14176
rect 4502 14112 4510 14176
rect 4190 13088 4510 14112
rect 4190 13024 4198 13088
rect 4262 13024 4278 13088
rect 4342 13024 4358 13088
rect 4422 13024 4438 13088
rect 4502 13024 4510 13088
rect 4190 12000 4510 13024
rect 4190 11936 4198 12000
rect 4262 11936 4278 12000
rect 4342 11936 4358 12000
rect 4422 11936 4438 12000
rect 4502 11936 4510 12000
rect 4190 10912 4510 11936
rect 4190 10848 4198 10912
rect 4262 10848 4278 10912
rect 4342 10848 4358 10912
rect 4422 10848 4438 10912
rect 4502 10848 4510 10912
rect 4190 9824 4510 10848
rect 4190 9760 4198 9824
rect 4262 9760 4278 9824
rect 4342 9760 4358 9824
rect 4422 9760 4438 9824
rect 4502 9760 4510 9824
rect 4190 8736 4510 9760
rect 4190 8672 4198 8736
rect 4262 8672 4278 8736
rect 4342 8672 4358 8736
rect 4422 8672 4438 8736
rect 4502 8672 4510 8736
rect 4190 7648 4510 8672
rect 4190 7584 4198 7648
rect 4262 7584 4278 7648
rect 4342 7584 4358 7648
rect 4422 7584 4438 7648
rect 4502 7584 4510 7648
rect 4190 6560 4510 7584
rect 4190 6496 4198 6560
rect 4262 6496 4278 6560
rect 4342 6496 4358 6560
rect 4422 6496 4438 6560
rect 4502 6496 4510 6560
rect 4190 5472 4510 6496
rect 4190 5408 4198 5472
rect 4262 5408 4278 5472
rect 4342 5408 4358 5472
rect 4422 5408 4438 5472
rect 4502 5408 4510 5472
rect 4190 4384 4510 5408
rect 4190 4320 4198 4384
rect 4262 4320 4278 4384
rect 4342 4320 4358 4384
rect 4422 4320 4438 4384
rect 4502 4320 4510 4384
rect 4190 3296 4510 4320
rect 4190 3232 4198 3296
rect 4262 3232 4278 3296
rect 4342 3232 4358 3296
rect 4422 3232 4438 3296
rect 4502 3232 4510 3296
rect 4190 2208 4510 3232
rect 4190 2144 4198 2208
rect 4262 2144 4278 2208
rect 4342 2144 4358 2208
rect 4422 2144 4438 2208
rect 4502 2144 4510 2208
rect 4190 2128 4510 2144
rect 19550 57152 19870 57712
rect 19550 57088 19558 57152
rect 19622 57088 19638 57152
rect 19702 57088 19718 57152
rect 19782 57088 19798 57152
rect 19862 57088 19870 57152
rect 19550 56064 19870 57088
rect 19550 56000 19558 56064
rect 19622 56000 19638 56064
rect 19702 56000 19718 56064
rect 19782 56000 19798 56064
rect 19862 56000 19870 56064
rect 19550 54976 19870 56000
rect 19550 54912 19558 54976
rect 19622 54912 19638 54976
rect 19702 54912 19718 54976
rect 19782 54912 19798 54976
rect 19862 54912 19870 54976
rect 19550 53888 19870 54912
rect 19550 53824 19558 53888
rect 19622 53824 19638 53888
rect 19702 53824 19718 53888
rect 19782 53824 19798 53888
rect 19862 53824 19870 53888
rect 19550 52800 19870 53824
rect 19550 52736 19558 52800
rect 19622 52736 19638 52800
rect 19702 52736 19718 52800
rect 19782 52736 19798 52800
rect 19862 52736 19870 52800
rect 19550 51712 19870 52736
rect 19550 51648 19558 51712
rect 19622 51648 19638 51712
rect 19702 51648 19718 51712
rect 19782 51648 19798 51712
rect 19862 51648 19870 51712
rect 19550 50624 19870 51648
rect 19550 50560 19558 50624
rect 19622 50560 19638 50624
rect 19702 50560 19718 50624
rect 19782 50560 19798 50624
rect 19862 50560 19870 50624
rect 19550 49536 19870 50560
rect 19550 49472 19558 49536
rect 19622 49472 19638 49536
rect 19702 49472 19718 49536
rect 19782 49472 19798 49536
rect 19862 49472 19870 49536
rect 19550 48448 19870 49472
rect 19550 48384 19558 48448
rect 19622 48384 19638 48448
rect 19702 48384 19718 48448
rect 19782 48384 19798 48448
rect 19862 48384 19870 48448
rect 19550 47360 19870 48384
rect 19550 47296 19558 47360
rect 19622 47296 19638 47360
rect 19702 47296 19718 47360
rect 19782 47296 19798 47360
rect 19862 47296 19870 47360
rect 19550 46272 19870 47296
rect 19550 46208 19558 46272
rect 19622 46208 19638 46272
rect 19702 46208 19718 46272
rect 19782 46208 19798 46272
rect 19862 46208 19870 46272
rect 19550 45184 19870 46208
rect 19550 45120 19558 45184
rect 19622 45120 19638 45184
rect 19702 45120 19718 45184
rect 19782 45120 19798 45184
rect 19862 45120 19870 45184
rect 19550 44096 19870 45120
rect 19550 44032 19558 44096
rect 19622 44032 19638 44096
rect 19702 44032 19718 44096
rect 19782 44032 19798 44096
rect 19862 44032 19870 44096
rect 19550 43008 19870 44032
rect 19550 42944 19558 43008
rect 19622 42944 19638 43008
rect 19702 42944 19718 43008
rect 19782 42944 19798 43008
rect 19862 42944 19870 43008
rect 19550 41920 19870 42944
rect 19550 41856 19558 41920
rect 19622 41856 19638 41920
rect 19702 41856 19718 41920
rect 19782 41856 19798 41920
rect 19862 41856 19870 41920
rect 19550 40832 19870 41856
rect 19550 40768 19558 40832
rect 19622 40768 19638 40832
rect 19702 40768 19718 40832
rect 19782 40768 19798 40832
rect 19862 40768 19870 40832
rect 19550 39744 19870 40768
rect 19550 39680 19558 39744
rect 19622 39680 19638 39744
rect 19702 39680 19718 39744
rect 19782 39680 19798 39744
rect 19862 39680 19870 39744
rect 19550 38656 19870 39680
rect 19550 38592 19558 38656
rect 19622 38592 19638 38656
rect 19702 38592 19718 38656
rect 19782 38592 19798 38656
rect 19862 38592 19870 38656
rect 19550 37568 19870 38592
rect 19550 37504 19558 37568
rect 19622 37504 19638 37568
rect 19702 37504 19718 37568
rect 19782 37504 19798 37568
rect 19862 37504 19870 37568
rect 19550 36480 19870 37504
rect 19550 36416 19558 36480
rect 19622 36416 19638 36480
rect 19702 36416 19718 36480
rect 19782 36416 19798 36480
rect 19862 36416 19870 36480
rect 19550 35392 19870 36416
rect 19550 35328 19558 35392
rect 19622 35328 19638 35392
rect 19702 35328 19718 35392
rect 19782 35328 19798 35392
rect 19862 35328 19870 35392
rect 19550 34304 19870 35328
rect 19550 34240 19558 34304
rect 19622 34240 19638 34304
rect 19702 34240 19718 34304
rect 19782 34240 19798 34304
rect 19862 34240 19870 34304
rect 19550 33216 19870 34240
rect 19550 33152 19558 33216
rect 19622 33152 19638 33216
rect 19702 33152 19718 33216
rect 19782 33152 19798 33216
rect 19862 33152 19870 33216
rect 19550 32128 19870 33152
rect 19550 32064 19558 32128
rect 19622 32064 19638 32128
rect 19702 32064 19718 32128
rect 19782 32064 19798 32128
rect 19862 32064 19870 32128
rect 19550 31040 19870 32064
rect 19550 30976 19558 31040
rect 19622 30976 19638 31040
rect 19702 30976 19718 31040
rect 19782 30976 19798 31040
rect 19862 30976 19870 31040
rect 19550 29952 19870 30976
rect 19550 29888 19558 29952
rect 19622 29888 19638 29952
rect 19702 29888 19718 29952
rect 19782 29888 19798 29952
rect 19862 29888 19870 29952
rect 19550 28864 19870 29888
rect 19550 28800 19558 28864
rect 19622 28800 19638 28864
rect 19702 28800 19718 28864
rect 19782 28800 19798 28864
rect 19862 28800 19870 28864
rect 19550 27776 19870 28800
rect 19550 27712 19558 27776
rect 19622 27712 19638 27776
rect 19702 27712 19718 27776
rect 19782 27712 19798 27776
rect 19862 27712 19870 27776
rect 19550 26688 19870 27712
rect 19550 26624 19558 26688
rect 19622 26624 19638 26688
rect 19702 26624 19718 26688
rect 19782 26624 19798 26688
rect 19862 26624 19870 26688
rect 19550 25600 19870 26624
rect 19550 25536 19558 25600
rect 19622 25536 19638 25600
rect 19702 25536 19718 25600
rect 19782 25536 19798 25600
rect 19862 25536 19870 25600
rect 19550 24512 19870 25536
rect 19550 24448 19558 24512
rect 19622 24448 19638 24512
rect 19702 24448 19718 24512
rect 19782 24448 19798 24512
rect 19862 24448 19870 24512
rect 19550 23424 19870 24448
rect 19550 23360 19558 23424
rect 19622 23360 19638 23424
rect 19702 23360 19718 23424
rect 19782 23360 19798 23424
rect 19862 23360 19870 23424
rect 19550 22336 19870 23360
rect 34910 57696 35230 57712
rect 34910 57632 34918 57696
rect 34982 57632 34998 57696
rect 35062 57632 35078 57696
rect 35142 57632 35158 57696
rect 35222 57632 35230 57696
rect 34910 56608 35230 57632
rect 34910 56544 34918 56608
rect 34982 56544 34998 56608
rect 35062 56544 35078 56608
rect 35142 56544 35158 56608
rect 35222 56544 35230 56608
rect 34910 55520 35230 56544
rect 34910 55456 34918 55520
rect 34982 55456 34998 55520
rect 35062 55456 35078 55520
rect 35142 55456 35158 55520
rect 35222 55456 35230 55520
rect 34910 54432 35230 55456
rect 34910 54368 34918 54432
rect 34982 54368 34998 54432
rect 35062 54368 35078 54432
rect 35142 54368 35158 54432
rect 35222 54368 35230 54432
rect 34910 53344 35230 54368
rect 34910 53280 34918 53344
rect 34982 53280 34998 53344
rect 35062 53280 35078 53344
rect 35142 53280 35158 53344
rect 35222 53280 35230 53344
rect 34910 52256 35230 53280
rect 34910 52192 34918 52256
rect 34982 52192 34998 52256
rect 35062 52192 35078 52256
rect 35142 52192 35158 52256
rect 35222 52192 35230 52256
rect 34910 51168 35230 52192
rect 34910 51104 34918 51168
rect 34982 51104 34998 51168
rect 35062 51104 35078 51168
rect 35142 51104 35158 51168
rect 35222 51104 35230 51168
rect 34910 50080 35230 51104
rect 34910 50016 34918 50080
rect 34982 50016 34998 50080
rect 35062 50016 35078 50080
rect 35142 50016 35158 50080
rect 35222 50016 35230 50080
rect 34910 48992 35230 50016
rect 34910 48928 34918 48992
rect 34982 48928 34998 48992
rect 35062 48928 35078 48992
rect 35142 48928 35158 48992
rect 35222 48928 35230 48992
rect 34910 47904 35230 48928
rect 34910 47840 34918 47904
rect 34982 47840 34998 47904
rect 35062 47840 35078 47904
rect 35142 47840 35158 47904
rect 35222 47840 35230 47904
rect 34910 46816 35230 47840
rect 34910 46752 34918 46816
rect 34982 46752 34998 46816
rect 35062 46752 35078 46816
rect 35142 46752 35158 46816
rect 35222 46752 35230 46816
rect 34910 45728 35230 46752
rect 34910 45664 34918 45728
rect 34982 45664 34998 45728
rect 35062 45664 35078 45728
rect 35142 45664 35158 45728
rect 35222 45664 35230 45728
rect 34910 44640 35230 45664
rect 34910 44576 34918 44640
rect 34982 44576 34998 44640
rect 35062 44576 35078 44640
rect 35142 44576 35158 44640
rect 35222 44576 35230 44640
rect 34910 43552 35230 44576
rect 50270 57152 50590 57712
rect 50270 57088 50278 57152
rect 50342 57088 50358 57152
rect 50422 57088 50438 57152
rect 50502 57088 50518 57152
rect 50582 57088 50590 57152
rect 50270 56064 50590 57088
rect 50270 56000 50278 56064
rect 50342 56000 50358 56064
rect 50422 56000 50438 56064
rect 50502 56000 50518 56064
rect 50582 56000 50590 56064
rect 50270 54976 50590 56000
rect 50270 54912 50278 54976
rect 50342 54912 50358 54976
rect 50422 54912 50438 54976
rect 50502 54912 50518 54976
rect 50582 54912 50590 54976
rect 50270 53888 50590 54912
rect 50270 53824 50278 53888
rect 50342 53824 50358 53888
rect 50422 53824 50438 53888
rect 50502 53824 50518 53888
rect 50582 53824 50590 53888
rect 50270 52800 50590 53824
rect 50270 52736 50278 52800
rect 50342 52736 50358 52800
rect 50422 52736 50438 52800
rect 50502 52736 50518 52800
rect 50582 52736 50590 52800
rect 50270 51712 50590 52736
rect 50270 51648 50278 51712
rect 50342 51648 50358 51712
rect 50422 51648 50438 51712
rect 50502 51648 50518 51712
rect 50582 51648 50590 51712
rect 50270 50624 50590 51648
rect 50270 50560 50278 50624
rect 50342 50560 50358 50624
rect 50422 50560 50438 50624
rect 50502 50560 50518 50624
rect 50582 50560 50590 50624
rect 50270 49536 50590 50560
rect 50270 49472 50278 49536
rect 50342 49472 50358 49536
rect 50422 49472 50438 49536
rect 50502 49472 50518 49536
rect 50582 49472 50590 49536
rect 50270 48448 50590 49472
rect 50270 48384 50278 48448
rect 50342 48384 50358 48448
rect 50422 48384 50438 48448
rect 50502 48384 50518 48448
rect 50582 48384 50590 48448
rect 50270 47360 50590 48384
rect 50270 47296 50278 47360
rect 50342 47296 50358 47360
rect 50422 47296 50438 47360
rect 50502 47296 50518 47360
rect 50582 47296 50590 47360
rect 50270 46272 50590 47296
rect 50270 46208 50278 46272
rect 50342 46208 50358 46272
rect 50422 46208 50438 46272
rect 50502 46208 50518 46272
rect 50582 46208 50590 46272
rect 50270 45184 50590 46208
rect 50270 45120 50278 45184
rect 50342 45120 50358 45184
rect 50422 45120 50438 45184
rect 50502 45120 50518 45184
rect 50582 45120 50590 45184
rect 38865 44164 38931 44165
rect 38865 44100 38866 44164
rect 38930 44100 38931 44164
rect 38865 44099 38931 44100
rect 34910 43488 34918 43552
rect 34982 43488 34998 43552
rect 35062 43488 35078 43552
rect 35142 43488 35158 43552
rect 35222 43488 35230 43552
rect 34910 42464 35230 43488
rect 34910 42400 34918 42464
rect 34982 42400 34998 42464
rect 35062 42400 35078 42464
rect 35142 42400 35158 42464
rect 35222 42400 35230 42464
rect 34910 41376 35230 42400
rect 34910 41312 34918 41376
rect 34982 41312 34998 41376
rect 35062 41312 35078 41376
rect 35142 41312 35158 41376
rect 35222 41312 35230 41376
rect 34910 40288 35230 41312
rect 34910 40224 34918 40288
rect 34982 40224 34998 40288
rect 35062 40224 35078 40288
rect 35142 40224 35158 40288
rect 35222 40224 35230 40288
rect 34910 39200 35230 40224
rect 34910 39136 34918 39200
rect 34982 39136 34998 39200
rect 35062 39136 35078 39200
rect 35142 39136 35158 39200
rect 35222 39136 35230 39200
rect 34910 38112 35230 39136
rect 34910 38048 34918 38112
rect 34982 38048 34998 38112
rect 35062 38048 35078 38112
rect 35142 38048 35158 38112
rect 35222 38048 35230 38112
rect 34910 37024 35230 38048
rect 34910 36960 34918 37024
rect 34982 36960 34998 37024
rect 35062 36960 35078 37024
rect 35142 36960 35158 37024
rect 35222 36960 35230 37024
rect 34910 35936 35230 36960
rect 34910 35872 34918 35936
rect 34982 35872 34998 35936
rect 35062 35872 35078 35936
rect 35142 35872 35158 35936
rect 35222 35872 35230 35936
rect 34910 34848 35230 35872
rect 34910 34784 34918 34848
rect 34982 34784 34998 34848
rect 35062 34784 35078 34848
rect 35142 34784 35158 34848
rect 35222 34784 35230 34848
rect 34910 33760 35230 34784
rect 34910 33696 34918 33760
rect 34982 33696 34998 33760
rect 35062 33696 35078 33760
rect 35142 33696 35158 33760
rect 35222 33696 35230 33760
rect 34910 32672 35230 33696
rect 34910 32608 34918 32672
rect 34982 32608 34998 32672
rect 35062 32608 35078 32672
rect 35142 32608 35158 32672
rect 35222 32608 35230 32672
rect 34910 31584 35230 32608
rect 34910 31520 34918 31584
rect 34982 31520 34998 31584
rect 35062 31520 35078 31584
rect 35142 31520 35158 31584
rect 35222 31520 35230 31584
rect 34910 30496 35230 31520
rect 34910 30432 34918 30496
rect 34982 30432 34998 30496
rect 35062 30432 35078 30496
rect 35142 30432 35158 30496
rect 35222 30432 35230 30496
rect 34910 29408 35230 30432
rect 34910 29344 34918 29408
rect 34982 29344 34998 29408
rect 35062 29344 35078 29408
rect 35142 29344 35158 29408
rect 35222 29344 35230 29408
rect 34910 28320 35230 29344
rect 34910 28256 34918 28320
rect 34982 28256 34998 28320
rect 35062 28256 35078 28320
rect 35142 28256 35158 28320
rect 35222 28256 35230 28320
rect 34910 27232 35230 28256
rect 34910 27168 34918 27232
rect 34982 27168 34998 27232
rect 35062 27168 35078 27232
rect 35142 27168 35158 27232
rect 35222 27168 35230 27232
rect 34910 26144 35230 27168
rect 38868 26349 38928 44099
rect 50270 44096 50590 45120
rect 50270 44032 50278 44096
rect 50342 44032 50358 44096
rect 50422 44032 50438 44096
rect 50502 44032 50518 44096
rect 50582 44032 50590 44096
rect 50270 43008 50590 44032
rect 50270 42944 50278 43008
rect 50342 42944 50358 43008
rect 50422 42944 50438 43008
rect 50502 42944 50518 43008
rect 50582 42944 50590 43008
rect 50270 41920 50590 42944
rect 50270 41856 50278 41920
rect 50342 41856 50358 41920
rect 50422 41856 50438 41920
rect 50502 41856 50518 41920
rect 50582 41856 50590 41920
rect 50270 40832 50590 41856
rect 50270 40768 50278 40832
rect 50342 40768 50358 40832
rect 50422 40768 50438 40832
rect 50502 40768 50518 40832
rect 50582 40768 50590 40832
rect 50270 39744 50590 40768
rect 50270 39680 50278 39744
rect 50342 39680 50358 39744
rect 50422 39680 50438 39744
rect 50502 39680 50518 39744
rect 50582 39680 50590 39744
rect 50270 38656 50590 39680
rect 50270 38592 50278 38656
rect 50342 38592 50358 38656
rect 50422 38592 50438 38656
rect 50502 38592 50518 38656
rect 50582 38592 50590 38656
rect 50270 37568 50590 38592
rect 50270 37504 50278 37568
rect 50342 37504 50358 37568
rect 50422 37504 50438 37568
rect 50502 37504 50518 37568
rect 50582 37504 50590 37568
rect 50270 36480 50590 37504
rect 50270 36416 50278 36480
rect 50342 36416 50358 36480
rect 50422 36416 50438 36480
rect 50502 36416 50518 36480
rect 50582 36416 50590 36480
rect 50270 35392 50590 36416
rect 50270 35328 50278 35392
rect 50342 35328 50358 35392
rect 50422 35328 50438 35392
rect 50502 35328 50518 35392
rect 50582 35328 50590 35392
rect 50270 34304 50590 35328
rect 50270 34240 50278 34304
rect 50342 34240 50358 34304
rect 50422 34240 50438 34304
rect 50502 34240 50518 34304
rect 50582 34240 50590 34304
rect 50270 33216 50590 34240
rect 50270 33152 50278 33216
rect 50342 33152 50358 33216
rect 50422 33152 50438 33216
rect 50502 33152 50518 33216
rect 50582 33152 50590 33216
rect 50270 32128 50590 33152
rect 50270 32064 50278 32128
rect 50342 32064 50358 32128
rect 50422 32064 50438 32128
rect 50502 32064 50518 32128
rect 50582 32064 50590 32128
rect 50270 31040 50590 32064
rect 50270 30976 50278 31040
rect 50342 30976 50358 31040
rect 50422 30976 50438 31040
rect 50502 30976 50518 31040
rect 50582 30976 50590 31040
rect 50270 29952 50590 30976
rect 50270 29888 50278 29952
rect 50342 29888 50358 29952
rect 50422 29888 50438 29952
rect 50502 29888 50518 29952
rect 50582 29888 50590 29952
rect 50270 28864 50590 29888
rect 50270 28800 50278 28864
rect 50342 28800 50358 28864
rect 50422 28800 50438 28864
rect 50502 28800 50518 28864
rect 50582 28800 50590 28864
rect 50270 27776 50590 28800
rect 50270 27712 50278 27776
rect 50342 27712 50358 27776
rect 50422 27712 50438 27776
rect 50502 27712 50518 27776
rect 50582 27712 50590 27776
rect 50270 26688 50590 27712
rect 50270 26624 50278 26688
rect 50342 26624 50358 26688
rect 50422 26624 50438 26688
rect 50502 26624 50518 26688
rect 50582 26624 50590 26688
rect 38865 26348 38931 26349
rect 38865 26284 38866 26348
rect 38930 26284 38931 26348
rect 38865 26283 38931 26284
rect 34910 26080 34918 26144
rect 34982 26080 34998 26144
rect 35062 26080 35078 26144
rect 35142 26080 35158 26144
rect 35222 26080 35230 26144
rect 34910 25056 35230 26080
rect 34910 24992 34918 25056
rect 34982 24992 34998 25056
rect 35062 24992 35078 25056
rect 35142 24992 35158 25056
rect 35222 24992 35230 25056
rect 34910 23968 35230 24992
rect 34910 23904 34918 23968
rect 34982 23904 34998 23968
rect 35062 23904 35078 23968
rect 35142 23904 35158 23968
rect 35222 23904 35230 23968
rect 23409 23356 23475 23357
rect 23409 23292 23410 23356
rect 23474 23292 23475 23356
rect 23409 23291 23475 23292
rect 19550 22272 19558 22336
rect 19622 22272 19638 22336
rect 19702 22272 19718 22336
rect 19782 22272 19798 22336
rect 19862 22272 19870 22336
rect 19550 21248 19870 22272
rect 19550 21184 19558 21248
rect 19622 21184 19638 21248
rect 19702 21184 19718 21248
rect 19782 21184 19798 21248
rect 19862 21184 19870 21248
rect 19550 20160 19870 21184
rect 19550 20096 19558 20160
rect 19622 20096 19638 20160
rect 19702 20096 19718 20160
rect 19782 20096 19798 20160
rect 19862 20096 19870 20160
rect 19550 19072 19870 20096
rect 19550 19008 19558 19072
rect 19622 19008 19638 19072
rect 19702 19008 19718 19072
rect 19782 19008 19798 19072
rect 19862 19008 19870 19072
rect 19550 17984 19870 19008
rect 19550 17920 19558 17984
rect 19622 17920 19638 17984
rect 19702 17920 19718 17984
rect 19782 17920 19798 17984
rect 19862 17920 19870 17984
rect 19550 16896 19870 17920
rect 19550 16832 19558 16896
rect 19622 16832 19638 16896
rect 19702 16832 19718 16896
rect 19782 16832 19798 16896
rect 19862 16832 19870 16896
rect 19550 15808 19870 16832
rect 19550 15744 19558 15808
rect 19622 15744 19638 15808
rect 19702 15744 19718 15808
rect 19782 15744 19798 15808
rect 19862 15744 19870 15808
rect 19550 14720 19870 15744
rect 23412 15197 23472 23291
rect 34910 22880 35230 23904
rect 34910 22816 34918 22880
rect 34982 22816 34998 22880
rect 35062 22816 35078 22880
rect 35142 22816 35158 22880
rect 35222 22816 35230 22880
rect 34910 21792 35230 22816
rect 34910 21728 34918 21792
rect 34982 21728 34998 21792
rect 35062 21728 35078 21792
rect 35142 21728 35158 21792
rect 35222 21728 35230 21792
rect 34910 20704 35230 21728
rect 34910 20640 34918 20704
rect 34982 20640 34998 20704
rect 35062 20640 35078 20704
rect 35142 20640 35158 20704
rect 35222 20640 35230 20704
rect 34910 19616 35230 20640
rect 34910 19552 34918 19616
rect 34982 19552 34998 19616
rect 35062 19552 35078 19616
rect 35142 19552 35158 19616
rect 35222 19552 35230 19616
rect 34910 18528 35230 19552
rect 34910 18464 34918 18528
rect 34982 18464 34998 18528
rect 35062 18464 35078 18528
rect 35142 18464 35158 18528
rect 35222 18464 35230 18528
rect 34910 17440 35230 18464
rect 34910 17376 34918 17440
rect 34982 17376 34998 17440
rect 35062 17376 35078 17440
rect 35142 17376 35158 17440
rect 35222 17376 35230 17440
rect 34910 16352 35230 17376
rect 34910 16288 34918 16352
rect 34982 16288 34998 16352
rect 35062 16288 35078 16352
rect 35142 16288 35158 16352
rect 35222 16288 35230 16352
rect 34910 15264 35230 16288
rect 34910 15200 34918 15264
rect 34982 15200 34998 15264
rect 35062 15200 35078 15264
rect 35142 15200 35158 15264
rect 35222 15200 35230 15264
rect 23409 15196 23475 15197
rect 23409 15132 23410 15196
rect 23474 15132 23475 15196
rect 23409 15131 23475 15132
rect 19550 14656 19558 14720
rect 19622 14656 19638 14720
rect 19702 14656 19718 14720
rect 19782 14656 19798 14720
rect 19862 14656 19870 14720
rect 19550 13632 19870 14656
rect 19550 13568 19558 13632
rect 19622 13568 19638 13632
rect 19702 13568 19718 13632
rect 19782 13568 19798 13632
rect 19862 13568 19870 13632
rect 19550 12544 19870 13568
rect 19550 12480 19558 12544
rect 19622 12480 19638 12544
rect 19702 12480 19718 12544
rect 19782 12480 19798 12544
rect 19862 12480 19870 12544
rect 19550 11456 19870 12480
rect 19550 11392 19558 11456
rect 19622 11392 19638 11456
rect 19702 11392 19718 11456
rect 19782 11392 19798 11456
rect 19862 11392 19870 11456
rect 19550 10368 19870 11392
rect 19550 10304 19558 10368
rect 19622 10304 19638 10368
rect 19702 10304 19718 10368
rect 19782 10304 19798 10368
rect 19862 10304 19870 10368
rect 19550 9280 19870 10304
rect 19550 9216 19558 9280
rect 19622 9216 19638 9280
rect 19702 9216 19718 9280
rect 19782 9216 19798 9280
rect 19862 9216 19870 9280
rect 19550 8192 19870 9216
rect 19550 8128 19558 8192
rect 19622 8128 19638 8192
rect 19702 8128 19718 8192
rect 19782 8128 19798 8192
rect 19862 8128 19870 8192
rect 19550 7104 19870 8128
rect 34910 14176 35230 15200
rect 34910 14112 34918 14176
rect 34982 14112 34998 14176
rect 35062 14112 35078 14176
rect 35142 14112 35158 14176
rect 35222 14112 35230 14176
rect 34910 13088 35230 14112
rect 34910 13024 34918 13088
rect 34982 13024 34998 13088
rect 35062 13024 35078 13088
rect 35142 13024 35158 13088
rect 35222 13024 35230 13088
rect 34910 12000 35230 13024
rect 34910 11936 34918 12000
rect 34982 11936 34998 12000
rect 35062 11936 35078 12000
rect 35142 11936 35158 12000
rect 35222 11936 35230 12000
rect 34910 10912 35230 11936
rect 34910 10848 34918 10912
rect 34982 10848 34998 10912
rect 35062 10848 35078 10912
rect 35142 10848 35158 10912
rect 35222 10848 35230 10912
rect 34910 9824 35230 10848
rect 34910 9760 34918 9824
rect 34982 9760 34998 9824
rect 35062 9760 35078 9824
rect 35142 9760 35158 9824
rect 35222 9760 35230 9824
rect 34910 8736 35230 9760
rect 34910 8672 34918 8736
rect 34982 8672 34998 8736
rect 35062 8672 35078 8736
rect 35142 8672 35158 8736
rect 35222 8672 35230 8736
rect 20281 7716 20347 7717
rect 20281 7652 20282 7716
rect 20346 7652 20347 7716
rect 20281 7651 20347 7652
rect 19550 7040 19558 7104
rect 19622 7040 19638 7104
rect 19702 7040 19718 7104
rect 19782 7040 19798 7104
rect 19862 7040 19870 7104
rect 19550 6016 19870 7040
rect 19550 5952 19558 6016
rect 19622 5952 19638 6016
rect 19702 5952 19718 6016
rect 19782 5952 19798 6016
rect 19862 5952 19870 6016
rect 19550 4928 19870 5952
rect 19550 4864 19558 4928
rect 19622 4864 19638 4928
rect 19702 4864 19718 4928
rect 19782 4864 19798 4928
rect 19862 4864 19870 4928
rect 19550 3840 19870 4864
rect 19550 3776 19558 3840
rect 19622 3776 19638 3840
rect 19702 3776 19718 3840
rect 19782 3776 19798 3840
rect 19862 3776 19870 3840
rect 19550 2752 19870 3776
rect 19550 2688 19558 2752
rect 19622 2688 19638 2752
rect 19702 2688 19718 2752
rect 19782 2688 19798 2752
rect 19862 2688 19870 2752
rect 19550 2128 19870 2688
rect 20284 917 20344 7651
rect 34910 7648 35230 8672
rect 34910 7584 34918 7648
rect 34982 7584 34998 7648
rect 35062 7584 35078 7648
rect 35142 7584 35158 7648
rect 35222 7584 35230 7648
rect 34910 6560 35230 7584
rect 34910 6496 34918 6560
rect 34982 6496 34998 6560
rect 35062 6496 35078 6560
rect 35142 6496 35158 6560
rect 35222 6496 35230 6560
rect 34910 5472 35230 6496
rect 34910 5408 34918 5472
rect 34982 5408 34998 5472
rect 35062 5408 35078 5472
rect 35142 5408 35158 5472
rect 35222 5408 35230 5472
rect 34910 4384 35230 5408
rect 34910 4320 34918 4384
rect 34982 4320 34998 4384
rect 35062 4320 35078 4384
rect 35142 4320 35158 4384
rect 35222 4320 35230 4384
rect 34910 3296 35230 4320
rect 50270 25600 50590 26624
rect 50270 25536 50278 25600
rect 50342 25536 50358 25600
rect 50422 25536 50438 25600
rect 50502 25536 50518 25600
rect 50582 25536 50590 25600
rect 50270 24512 50590 25536
rect 50270 24448 50278 24512
rect 50342 24448 50358 24512
rect 50422 24448 50438 24512
rect 50502 24448 50518 24512
rect 50582 24448 50590 24512
rect 50270 23424 50590 24448
rect 50270 23360 50278 23424
rect 50342 23360 50358 23424
rect 50422 23360 50438 23424
rect 50502 23360 50518 23424
rect 50582 23360 50590 23424
rect 50270 22336 50590 23360
rect 50270 22272 50278 22336
rect 50342 22272 50358 22336
rect 50422 22272 50438 22336
rect 50502 22272 50518 22336
rect 50582 22272 50590 22336
rect 50270 21248 50590 22272
rect 50270 21184 50278 21248
rect 50342 21184 50358 21248
rect 50422 21184 50438 21248
rect 50502 21184 50518 21248
rect 50582 21184 50590 21248
rect 50270 20160 50590 21184
rect 50270 20096 50278 20160
rect 50342 20096 50358 20160
rect 50422 20096 50438 20160
rect 50502 20096 50518 20160
rect 50582 20096 50590 20160
rect 50270 19072 50590 20096
rect 50270 19008 50278 19072
rect 50342 19008 50358 19072
rect 50422 19008 50438 19072
rect 50502 19008 50518 19072
rect 50582 19008 50590 19072
rect 50270 17984 50590 19008
rect 50270 17920 50278 17984
rect 50342 17920 50358 17984
rect 50422 17920 50438 17984
rect 50502 17920 50518 17984
rect 50582 17920 50590 17984
rect 50270 16896 50590 17920
rect 50270 16832 50278 16896
rect 50342 16832 50358 16896
rect 50422 16832 50438 16896
rect 50502 16832 50518 16896
rect 50582 16832 50590 16896
rect 50270 15808 50590 16832
rect 50270 15744 50278 15808
rect 50342 15744 50358 15808
rect 50422 15744 50438 15808
rect 50502 15744 50518 15808
rect 50582 15744 50590 15808
rect 50270 14720 50590 15744
rect 50270 14656 50278 14720
rect 50342 14656 50358 14720
rect 50422 14656 50438 14720
rect 50502 14656 50518 14720
rect 50582 14656 50590 14720
rect 50270 13632 50590 14656
rect 50270 13568 50278 13632
rect 50342 13568 50358 13632
rect 50422 13568 50438 13632
rect 50502 13568 50518 13632
rect 50582 13568 50590 13632
rect 50270 12544 50590 13568
rect 50270 12480 50278 12544
rect 50342 12480 50358 12544
rect 50422 12480 50438 12544
rect 50502 12480 50518 12544
rect 50582 12480 50590 12544
rect 50270 11456 50590 12480
rect 50270 11392 50278 11456
rect 50342 11392 50358 11456
rect 50422 11392 50438 11456
rect 50502 11392 50518 11456
rect 50582 11392 50590 11456
rect 50270 10368 50590 11392
rect 50270 10304 50278 10368
rect 50342 10304 50358 10368
rect 50422 10304 50438 10368
rect 50502 10304 50518 10368
rect 50582 10304 50590 10368
rect 50270 9280 50590 10304
rect 50270 9216 50278 9280
rect 50342 9216 50358 9280
rect 50422 9216 50438 9280
rect 50502 9216 50518 9280
rect 50582 9216 50590 9280
rect 50270 8192 50590 9216
rect 50270 8128 50278 8192
rect 50342 8128 50358 8192
rect 50422 8128 50438 8192
rect 50502 8128 50518 8192
rect 50582 8128 50590 8192
rect 50270 7104 50590 8128
rect 50270 7040 50278 7104
rect 50342 7040 50358 7104
rect 50422 7040 50438 7104
rect 50502 7040 50518 7104
rect 50582 7040 50590 7104
rect 50270 6016 50590 7040
rect 50270 5952 50278 6016
rect 50342 5952 50358 6016
rect 50422 5952 50438 6016
rect 50502 5952 50518 6016
rect 50582 5952 50590 6016
rect 50270 4928 50590 5952
rect 50270 4864 50278 4928
rect 50342 4864 50358 4928
rect 50422 4864 50438 4928
rect 50502 4864 50518 4928
rect 50582 4864 50590 4928
rect 41257 3908 41323 3909
rect 41257 3844 41258 3908
rect 41322 3844 41323 3908
rect 41257 3843 41323 3844
rect 34910 3232 34918 3296
rect 34982 3232 34998 3296
rect 35062 3232 35078 3296
rect 35142 3232 35158 3296
rect 35222 3232 35230 3296
rect 34910 2208 35230 3232
rect 41260 2957 41320 3843
rect 50270 3840 50590 4864
rect 50270 3776 50278 3840
rect 50342 3776 50358 3840
rect 50422 3776 50438 3840
rect 50502 3776 50518 3840
rect 50582 3776 50590 3840
rect 41257 2956 41323 2957
rect 41257 2892 41258 2956
rect 41322 2892 41323 2956
rect 41257 2891 41323 2892
rect 34910 2144 34918 2208
rect 34982 2144 34998 2208
rect 35062 2144 35078 2208
rect 35142 2144 35158 2208
rect 35222 2144 35230 2208
rect 34910 2128 35230 2144
rect 50270 2752 50590 3776
rect 50270 2688 50278 2752
rect 50342 2688 50358 2752
rect 50422 2688 50438 2752
rect 50502 2688 50518 2752
rect 50582 2688 50590 2752
rect 50270 2128 50590 2688
rect 20281 916 20347 917
rect 20281 852 20282 916
rect 20346 852 20347 916
rect 20281 851 20347 852
use sky130_fd_sc_hd__decap_12  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 2466 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1607639953
transform 1 0 1362 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1607639953
transform 1 0 2466 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1607639953
transform 1 0 1362 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 1086 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1607639953
transform 1 0 1086 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1607639953
transform 1 0 4674 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1607639953
transform 1 0 3570 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1607639953
transform 1 0 5134 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1607639953
transform 1 0 4030 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 3570 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 3938 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1607639953
transform 1 0 6790 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 6514 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 5778 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp 1607639953
transform 1 0 6882 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 6238 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1607639953
transform 1 0 6698 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1607639953
transform 1 0 6790 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _203_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 7158 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_84
timestamp 1607639953
transform 1 0 8814 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_74
timestamp 1607639953
transform 1 0 7894 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_81
timestamp 1607639953
transform 1 0 8538 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1607639953
transform 1 0 7434 0 -1 2720
box -38 -48 1142 592
use AND2X1  AND2X1
timestamp 1608122862
transform 1 0 8078 0 1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_1_108
timestamp 1607639953
transform 1 0 11022 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_96
timestamp 1607639953
transform 1 0 9918 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1607639953
transform 1 0 10838 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1607639953
transform 1 0 9734 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1607639953
transform 1 0 9642 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1607639953
transform 1 0 12402 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1607639953
transform 1 0 12126 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1607639953
transform 1 0 12586 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1607639953
transform 1 0 11942 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1607639953
transform 1 0 12310 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1607639953
transform 1 0 12494 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1607639953
transform 1 0 14610 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1607639953
transform 1 0 13506 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1607639953
transform 1 0 14794 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1607639953
transform 1 0 13690 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1607639953
transform 1 0 16818 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1607639953
transform 1 0 15714 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1607639953
transform 1 0 16542 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1607639953
transform 1 0 15438 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1607639953
transform 1 0 15346 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_191
timestamp 1607639953
transform 1 0 18658 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_184
timestamp 1607639953
transform 1 0 18014 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_195
timestamp 1607639953
transform 1 0 19026 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_187
timestamp 1607639953
transform 1 0 18290 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1607639953
transform 1 0 17646 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1607639953
transform 1 0 17922 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1607639953
transform 1 0 18198 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _167_
timestamp 1607639953
transform 1 0 19210 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1607639953
transform 1 0 18382 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_215
timestamp 1607639953
transform 1 0 20866 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_203
timestamp 1607639953
transform 1 0 19762 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1607639953
transform 1 0 21142 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_216 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 20958 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1607639953
transform 1 0 20590 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_200
timestamp 1607639953
transform 1 0 19486 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1607639953
transform 1 0 21050 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_239
timestamp 1607639953
transform 1 0 23074 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_227
timestamp 1607639953
transform 1 0 21970 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1607639953
transform 1 0 23350 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1607639953
transform 1 0 22246 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1607639953
transform 1 0 24730 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1607639953
transform 1 0 23626 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1607639953
transform 1 0 23442 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1607639953
transform 1 0 25098 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1607639953
transform 1 0 23994 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1607639953
transform 1 0 23534 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1607639953
transform 1 0 23902 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1607639953
transform 1 0 26938 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_269
timestamp 1607639953
transform 1 0 25834 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_280
timestamp 1607639953
transform 1 0 26846 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1607639953
transform 1 0 26202 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1607639953
transform 1 0 26754 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_306
timestamp 1607639953
transform 1 0 29238 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1607639953
transform 1 0 28042 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_304
timestamp 1607639953
transform 1 0 29054 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_292
timestamp 1607639953
transform 1 0 27950 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1607639953
transform 1 0 29146 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_330
timestamp 1607639953
transform 1 0 31446 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_318
timestamp 1607639953
transform 1 0 30342 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_323
timestamp 1607639953
transform 1 0 30802 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_311
timestamp 1607639953
transform 1 0 29698 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1607639953
transform 1 0 29606 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_342
timestamp 1607639953
transform 1 0 32550 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_342
timestamp 1607639953
transform 1 0 32550 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_335
timestamp 1607639953
transform 1 0 31906 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1607639953
transform 1 0 32458 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_367
timestamp 1607639953
transform 1 0 34850 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_354
timestamp 1607639953
transform 1 0 33654 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_373
timestamp 1607639953
transform 1 0 35402 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_366
timestamp 1607639953
transform 1 0 34758 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_354
timestamp 1607639953
transform 1 0 33654 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1607639953
transform 1 0 34758 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1607639953
transform 1 0 35310 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_391
timestamp 1607639953
transform 1 0 37058 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1607639953
transform 1 0 35954 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_385
timestamp 1607639953
transform 1 0 36506 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_415
timestamp 1607639953
transform 1 0 39266 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_403
timestamp 1607639953
transform 1 0 38162 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_416
timestamp 1607639953
transform 1 0 39358 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_404
timestamp 1607639953
transform 1 0 38254 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_397
timestamp 1607639953
transform 1 0 37610 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1607639953
transform 1 0 38162 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_440
timestamp 1607639953
transform 1 0 41566 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_428
timestamp 1607639953
transform 1 0 40462 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_435
timestamp 1607639953
transform 1 0 41106 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_428
timestamp 1607639953
transform 1 0 40462 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1607639953
transform 1 0 40370 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1607639953
transform 1 0 41014 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_452
timestamp 1607639953
transform 1 0 42670 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_459
timestamp 1607639953
transform 1 0 43314 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_447
timestamp 1607639953
transform 1 0 42210 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_476
timestamp 1607639953
transform 1 0 44878 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_464
timestamp 1607639953
transform 1 0 43774 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_478
timestamp 1607639953
transform 1 0 45062 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_466
timestamp 1607639953
transform 1 0 43958 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1607639953
transform 1 0 43866 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_501
timestamp 1607639953
transform 1 0 47178 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_489
timestamp 1607639953
transform 1 0 46074 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_497
timestamp 1607639953
transform 1 0 46810 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_490
timestamp 1607639953
transform 1 0 46166 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1607639953
transform 1 0 45982 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1607639953
transform 1 0 46718 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_525
timestamp 1607639953
transform 1 0 49386 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_513
timestamp 1607639953
transform 1 0 48282 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_528
timestamp 1607639953
transform 1 0 49662 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_521
timestamp 1607639953
transform 1 0 49018 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_509
timestamp 1607639953
transform 1 0 47914 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1607639953
transform 1 0 49570 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_550
timestamp 1607639953
transform 1 0 51686 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_537
timestamp 1607639953
transform 1 0 50490 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_546
timestamp 1607639953
transform 1 0 51318 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_534
timestamp 1607639953
transform 1 0 50214 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1607639953
transform 1 0 51594 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1607639953
transform 1 0 49938 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_562
timestamp 1607639953
transform 1 0 52790 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_571
timestamp 1607639953
transform 1 0 53618 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_559
timestamp 1607639953
transform 1 0 52514 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1607639953
transform 1 0 52422 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_586
timestamp 1607639953
transform 1 0 54998 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_574
timestamp 1607639953
transform 1 0 53894 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_590
timestamp 1607639953
transform 1 0 55366 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_583
timestamp 1607639953
transform 1 0 54722 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1607639953
transform 1 0 55274 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_611
timestamp 1607639953
transform 1 0 57298 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_598
timestamp 1607639953
transform 1 0 56102 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_614
timestamp 1607639953
transform 1 0 57574 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_602
timestamp 1607639953
transform 1 0 56470 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1607639953
transform 1 0 57206 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_623
timestamp 1607639953
transform 1 0 58402 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_621
timestamp 1607639953
transform 1 0 58218 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1607639953
transform 1 0 58126 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1607639953
transform -1 0 58862 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1607639953
transform -1 0 58862 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1607639953
transform 1 0 2466 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1607639953
transform 1 0 1362 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1607639953
transform 1 0 1086 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1607639953
transform 1 0 5134 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1607639953
transform 1 0 4030 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1607639953
transform 1 0 3570 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1607639953
transform 1 0 3938 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1607639953
transform 1 0 6238 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1607639953
transform 1 0 8446 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1607639953
transform 1 0 7342 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1607639953
transform 1 0 10746 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1607639953
transform 1 0 9642 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1607639953
transform 1 0 9550 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1607639953
transform 1 0 12954 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1607639953
transform 1 0 11850 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1607639953
transform 1 0 15254 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1607639953
transform 1 0 14058 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1607639953
transform 1 0 15162 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1607639953
transform 1 0 16358 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1607639953
transform 1 0 18566 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1607639953
transform 1 0 17462 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1607639953
transform 1 0 20866 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1607639953
transform 1 0 19670 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1607639953
transform 1 0 20774 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1607639953
transform 1 0 23074 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1607639953
transform 1 0 21970 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1607639953
transform 1 0 25282 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1607639953
transform 1 0 24178 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_276
timestamp 1607639953
transform 1 0 26478 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1607639953
transform 1 0 26386 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_300
timestamp 1607639953
transform 1 0 28686 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_288
timestamp 1607639953
transform 1 0 27582 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_324
timestamp 1607639953
transform 1 0 30894 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_312
timestamp 1607639953
transform 1 0 29790 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_349
timestamp 1607639953
transform 1 0 33194 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_337
timestamp 1607639953
transform 1 0 32090 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1607639953
transform 1 0 31998 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_373
timestamp 1607639953
transform 1 0 35402 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_361
timestamp 1607639953
transform 1 0 34298 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_385
timestamp 1607639953
transform 1 0 36506 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_410
timestamp 1607639953
transform 1 0 38806 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_398
timestamp 1607639953
transform 1 0 37702 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1607639953
transform 1 0 37610 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_434
timestamp 1607639953
transform 1 0 41014 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_422
timestamp 1607639953
transform 1 0 39910 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_459
timestamp 1607639953
transform 1 0 43314 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_446
timestamp 1607639953
transform 1 0 42118 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1607639953
transform 1 0 43222 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_483
timestamp 1607639953
transform 1 0 45522 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_471
timestamp 1607639953
transform 1 0 44418 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_495
timestamp 1607639953
transform 1 0 46626 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_520
timestamp 1607639953
transform 1 0 48926 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_507
timestamp 1607639953
transform 1 0 47730 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1607639953
transform 1 0 48834 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_544
timestamp 1607639953
transform 1 0 51134 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_532
timestamp 1607639953
transform 1 0 50030 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_570
timestamp 1607639953
transform 1 0 53526 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_558
timestamp 1607639953
transform 1 0 52422 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_552
timestamp 1607639953
transform 1 0 51870 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _139_
timestamp 1607639953
transform 1 0 52146 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_593
timestamp 1607639953
transform 1 0 55642 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_581
timestamp 1607639953
transform 1 0 54538 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_578
timestamp 1607639953
transform 1 0 54262 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1607639953
transform 1 0 54446 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_605
timestamp 1607639953
transform 1 0 56746 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_624
timestamp 1607639953
transform 1 0 58494 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_617
timestamp 1607639953
transform 1 0 57850 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1607639953
transform -1 0 58862 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _160_
timestamp 1607639953
transform 1 0 58218 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1607639953
transform 1 0 2466 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1607639953
transform 1 0 1362 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1607639953
transform 1 0 1086 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1607639953
transform 1 0 4674 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1607639953
transform 1 0 3570 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_66
timestamp 1607639953
transform 1 0 7158 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1607639953
transform 1 0 6790 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1607639953
transform 1 0 6514 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1607639953
transform 1 0 5778 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1607639953
transform 1 0 6698 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_84
timestamp 1607639953
transform 1 0 8814 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_70
timestamp 1607639953
transform 1 0 7526 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _100_
timestamp 1607639953
transform 1 0 7250 0 1 3808
box -38 -48 314 592
use AND2X2  AND2X2
timestamp 1608122862
transform 1 0 8078 0 1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_3_108
timestamp 1607639953
transform 1 0 11022 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_96
timestamp 1607639953
transform 1 0 9918 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1607639953
transform 1 0 12402 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1607639953
transform 1 0 12126 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1607639953
transform 1 0 12310 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1607639953
transform 1 0 14610 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1607639953
transform 1 0 13506 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1607639953
transform 1 0 16818 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1607639953
transform 1 0 15714 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1607639953
transform 1 0 19118 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1607639953
transform 1 0 18014 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1607639953
transform 1 0 17922 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1607639953
transform 1 0 21326 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1607639953
transform 1 0 20222 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1607639953
transform 1 0 22430 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1607639953
transform 1 0 24730 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1607639953
transform 1 0 23626 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1607639953
transform 1 0 23534 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1607639953
transform 1 0 26938 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_269
timestamp 1607639953
transform 1 0 25834 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_306
timestamp 1607639953
transform 1 0 29238 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1607639953
transform 1 0 28042 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1607639953
transform 1 0 29146 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_330
timestamp 1607639953
transform 1 0 31446 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_318
timestamp 1607639953
transform 1 0 30342 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_342
timestamp 1607639953
transform 1 0 32550 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_367
timestamp 1607639953
transform 1 0 34850 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_354
timestamp 1607639953
transform 1 0 33654 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1607639953
transform 1 0 34758 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_391
timestamp 1607639953
transform 1 0 37058 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_379
timestamp 1607639953
transform 1 0 35954 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_415
timestamp 1607639953
transform 1 0 39266 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_403
timestamp 1607639953
transform 1 0 38162 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_440
timestamp 1607639953
transform 1 0 41566 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_428
timestamp 1607639953
transform 1 0 40462 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1607639953
transform 1 0 40370 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_452
timestamp 1607639953
transform 1 0 42670 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_476
timestamp 1607639953
transform 1 0 44878 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_464
timestamp 1607639953
transform 1 0 43774 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_501
timestamp 1607639953
transform 1 0 47178 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_489
timestamp 1607639953
transform 1 0 46074 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1607639953
transform 1 0 45982 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_525
timestamp 1607639953
transform 1 0 49386 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_513
timestamp 1607639953
transform 1 0 48282 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_550
timestamp 1607639953
transform 1 0 51686 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_537
timestamp 1607639953
transform 1 0 50490 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1607639953
transform 1 0 51594 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_562
timestamp 1607639953
transform 1 0 52790 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_586
timestamp 1607639953
transform 1 0 54998 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_574
timestamp 1607639953
transform 1 0 53894 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_611
timestamp 1607639953
transform 1 0 57298 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_598
timestamp 1607639953
transform 1 0 56102 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1607639953
transform 1 0 57206 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_623
timestamp 1607639953
transform 1 0 58402 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1607639953
transform -1 0 58862 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1607639953
transform 1 0 2466 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1607639953
transform 1 0 1362 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1607639953
transform 1 0 1086 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1607639953
transform 1 0 5134 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1607639953
transform 1 0 4030 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1607639953
transform 1 0 3570 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1607639953
transform 1 0 3938 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1607639953
transform 1 0 6238 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1607639953
transform 1 0 8446 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1607639953
transform 1 0 7342 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1607639953
transform 1 0 10746 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1607639953
transform 1 0 9642 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1607639953
transform 1 0 9550 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1607639953
transform 1 0 12954 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1607639953
transform 1 0 11850 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1607639953
transform 1 0 15254 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1607639953
transform 1 0 14058 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1607639953
transform 1 0 15162 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1607639953
transform 1 0 16358 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1607639953
transform 1 0 18566 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1607639953
transform 1 0 17462 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1607639953
transform 1 0 20866 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1607639953
transform 1 0 19670 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1607639953
transform 1 0 20774 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1607639953
transform 1 0 23074 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1607639953
transform 1 0 21970 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1607639953
transform 1 0 25282 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1607639953
transform 1 0 24178 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_276
timestamp 1607639953
transform 1 0 26478 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1607639953
transform 1 0 26386 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_300
timestamp 1607639953
transform 1 0 28686 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_288
timestamp 1607639953
transform 1 0 27582 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_324
timestamp 1607639953
transform 1 0 30894 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_312
timestamp 1607639953
transform 1 0 29790 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_349
timestamp 1607639953
transform 1 0 33194 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_337
timestamp 1607639953
transform 1 0 32090 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1607639953
transform 1 0 31998 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_373
timestamp 1607639953
transform 1 0 35402 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_361
timestamp 1607639953
transform 1 0 34298 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_385
timestamp 1607639953
transform 1 0 36506 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_410
timestamp 1607639953
transform 1 0 38806 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_398
timestamp 1607639953
transform 1 0 37702 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1607639953
transform 1 0 37610 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_434
timestamp 1607639953
transform 1 0 41014 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_422
timestamp 1607639953
transform 1 0 39910 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_459
timestamp 1607639953
transform 1 0 43314 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_446
timestamp 1607639953
transform 1 0 42118 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1607639953
transform 1 0 43222 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_483
timestamp 1607639953
transform 1 0 45522 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_471
timestamp 1607639953
transform 1 0 44418 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_503
timestamp 1607639953
transform 1 0 47362 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_495
timestamp 1607639953
transform 1 0 46626 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _114_
timestamp 1607639953
transform 1 0 47454 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_520
timestamp 1607639953
transform 1 0 48926 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_507
timestamp 1607639953
transform 1 0 47730 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1607639953
transform 1 0 48834 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_544
timestamp 1607639953
transform 1 0 51134 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_532
timestamp 1607639953
transform 1 0 50030 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_568
timestamp 1607639953
transform 1 0 53342 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_556
timestamp 1607639953
transform 1 0 52238 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_593
timestamp 1607639953
transform 1 0 55642 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_581
timestamp 1607639953
transform 1 0 54538 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1607639953
transform 1 0 54446 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_605
timestamp 1607639953
transform 1 0 56746 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_617
timestamp 1607639953
transform 1 0 57850 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1607639953
transform -1 0 58862 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1607639953
transform 1 0 2466 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1607639953
transform 1 0 1362 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1607639953
transform 1 0 1086 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1607639953
transform 1 0 4674 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1607639953
transform 1 0 3570 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1607639953
transform 1 0 6790 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1607639953
transform 1 0 6514 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1607639953
transform 1 0 5778 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1607639953
transform 1 0 6698 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_84
timestamp 1607639953
transform 1 0 8814 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_74
timestamp 1607639953
transform 1 0 7894 0 1 4896
box -38 -48 222 592
use AOI21X1  AOI21X1
timestamp 1608122862
transform 1 0 8078 0 1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_5_108
timestamp 1607639953
transform 1 0 11022 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_96
timestamp 1607639953
transform 1 0 9918 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1607639953
transform 1 0 12402 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1607639953
transform 1 0 12126 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1607639953
transform 1 0 12310 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1607639953
transform 1 0 14610 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1607639953
transform 1 0 13506 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1607639953
transform 1 0 16818 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1607639953
transform 1 0 15714 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1607639953
transform 1 0 19118 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1607639953
transform 1 0 18014 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1607639953
transform 1 0 17922 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1607639953
transform 1 0 21326 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1607639953
transform 1 0 20222 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1607639953
transform 1 0 22430 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1607639953
transform 1 0 24730 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1607639953
transform 1 0 23626 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1607639953
transform 1 0 23534 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1607639953
transform 1 0 26938 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_269
timestamp 1607639953
transform 1 0 25834 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_306
timestamp 1607639953
transform 1 0 29238 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1607639953
transform 1 0 28042 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1607639953
transform 1 0 29146 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_330
timestamp 1607639953
transform 1 0 31446 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_318
timestamp 1607639953
transform 1 0 30342 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_342
timestamp 1607639953
transform 1 0 32550 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_367
timestamp 1607639953
transform 1 0 34850 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_354
timestamp 1607639953
transform 1 0 33654 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1607639953
transform 1 0 34758 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_391
timestamp 1607639953
transform 1 0 37058 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_379
timestamp 1607639953
transform 1 0 35954 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_415
timestamp 1607639953
transform 1 0 39266 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_403
timestamp 1607639953
transform 1 0 38162 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_440
timestamp 1607639953
transform 1 0 41566 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_428
timestamp 1607639953
transform 1 0 40462 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1607639953
transform 1 0 40370 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_452
timestamp 1607639953
transform 1 0 42670 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_476
timestamp 1607639953
transform 1 0 44878 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_464
timestamp 1607639953
transform 1 0 43774 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_501
timestamp 1607639953
transform 1 0 47178 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_489
timestamp 1607639953
transform 1 0 46074 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1607639953
transform 1 0 45982 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_525
timestamp 1607639953
transform 1 0 49386 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_513
timestamp 1607639953
transform 1 0 48282 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_550
timestamp 1607639953
transform 1 0 51686 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_537
timestamp 1607639953
transform 1 0 50490 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1607639953
transform 1 0 51594 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_562
timestamp 1607639953
transform 1 0 52790 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_586
timestamp 1607639953
transform 1 0 54998 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_574
timestamp 1607639953
transform 1 0 53894 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_611
timestamp 1607639953
transform 1 0 57298 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_598
timestamp 1607639953
transform 1 0 56102 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1607639953
transform 1 0 57206 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_623
timestamp 1607639953
transform 1 0 58402 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1607639953
transform -1 0 58862 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1607639953
transform 1 0 2466 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1607639953
transform 1 0 1362 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1607639953
transform 1 0 2466 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1607639953
transform 1 0 1362 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1607639953
transform 1 0 1086 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1607639953
transform 1 0 1086 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1607639953
transform 1 0 4674 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1607639953
transform 1 0 3570 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1607639953
transform 1 0 5134 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1607639953
transform 1 0 4030 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1607639953
transform 1 0 3570 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1607639953
transform 1 0 3938 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1607639953
transform 1 0 6790 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1607639953
transform 1 0 6514 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1607639953
transform 1 0 5778 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1607639953
transform 1 0 6238 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1607639953
transform 1 0 6698 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1607639953
transform 1 0 8998 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_74
timestamp 1607639953
transform 1 0 7894 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1607639953
transform 1 0 8446 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1607639953
transform 1 0 7342 0 -1 5984
box -38 -48 1142 592
use AOI22X1  AOI22X1
timestamp 1608122862
transform 1 0 8078 0 1 5984
box 0 -48 920 592
use sky130_fd_sc_hd__decap_12  FILLER_7_102
timestamp 1607639953
transform 1 0 10470 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_98
timestamp 1607639953
transform 1 0 10102 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1607639953
transform 1 0 10746 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1607639953
transform 1 0 9642 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1607639953
transform 1 0 9550 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _092_
timestamp 1607639953
transform 1 0 10194 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1607639953
transform 1 0 12402 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_114
timestamp 1607639953
transform 1 0 11574 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1607639953
transform 1 0 12954 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1607639953
transform 1 0 11850 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1607639953
transform 1 0 12310 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1607639953
transform 1 0 14610 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1607639953
transform 1 0 13506 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1607639953
transform 1 0 15254 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1607639953
transform 1 0 14058 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1607639953
transform 1 0 15162 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1607639953
transform 1 0 16818 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1607639953
transform 1 0 15714 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1607639953
transform 1 0 16358 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1607639953
transform 1 0 19118 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1607639953
transform 1 0 18014 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_195
timestamp 1607639953
transform 1 0 19026 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_190
timestamp 1607639953
transform 1 0 18566 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1607639953
transform 1 0 17462 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1607639953
transform 1 0 17922 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1607639953
transform 1 0 18750 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1607639953
transform 1 0 21326 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1607639953
transform 1 0 20222 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1607639953
transform 1 0 20866 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1607639953
transform 1 0 20682 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_207
timestamp 1607639953
transform 1 0 20130 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1607639953
transform 1 0 20774 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1607639953
transform 1 0 22430 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1607639953
transform 1 0 23074 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1607639953
transform 1 0 21970 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1607639953
transform 1 0 24730 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1607639953
transform 1 0 23626 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1607639953
transform 1 0 25282 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1607639953
transform 1 0 24178 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1607639953
transform 1 0 23534 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1607639953
transform 1 0 26938 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_269
timestamp 1607639953
transform 1 0 25834 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_276
timestamp 1607639953
transform 1 0 26478 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1607639953
transform 1 0 26386 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_306
timestamp 1607639953
transform 1 0 29238 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1607639953
transform 1 0 28042 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_299
timestamp 1607639953
transform 1 0 28594 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_288
timestamp 1607639953
transform 1 0 27582 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1607639953
transform 1 0 29146 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _000_
timestamp 1607639953
transform 1 0 28318 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_330
timestamp 1607639953
transform 1 0 31446 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_318
timestamp 1607639953
transform 1 0 30342 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_323
timestamp 1607639953
transform 1 0 30802 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_311
timestamp 1607639953
transform 1 0 29698 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_342
timestamp 1607639953
transform 1 0 32550 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_349
timestamp 1607639953
transform 1 0 33194 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_337
timestamp 1607639953
transform 1 0 32090 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_335
timestamp 1607639953
transform 1 0 31906 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1607639953
transform 1 0 31998 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_367
timestamp 1607639953
transform 1 0 34850 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_354
timestamp 1607639953
transform 1 0 33654 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_373
timestamp 1607639953
transform 1 0 35402 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_361
timestamp 1607639953
transform 1 0 34298 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1607639953
transform 1 0 34758 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_386
timestamp 1607639953
transform 1 0 36598 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_379
timestamp 1607639953
transform 1 0 35954 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_385
timestamp 1607639953
transform 1 0 36506 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _199_
timestamp 1607639953
transform 1 0 36322 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_410
timestamp 1607639953
transform 1 0 38806 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_398
timestamp 1607639953
transform 1 0 37702 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_410
timestamp 1607639953
transform 1 0 38806 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_398
timestamp 1607639953
transform 1 0 37702 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1607639953
transform 1 0 37610 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_440
timestamp 1607639953
transform 1 0 41566 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_428
timestamp 1607639953
transform 1 0 40462 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_426
timestamp 1607639953
transform 1 0 40278 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_422
timestamp 1607639953
transform 1 0 39910 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_434
timestamp 1607639953
transform 1 0 41014 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_422
timestamp 1607639953
transform 1 0 39910 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1607639953
transform 1 0 40370 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_452
timestamp 1607639953
transform 1 0 42670 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_462
timestamp 1607639953
transform 1 0 43590 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_446
timestamp 1607639953
transform 1 0 42118 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1607639953
transform 1 0 43222 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _182_
timestamp 1607639953
transform 1 0 43314 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_476
timestamp 1607639953
transform 1 0 44878 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_464
timestamp 1607639953
transform 1 0 43774 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_474
timestamp 1607639953
transform 1 0 44694 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_501
timestamp 1607639953
transform 1 0 47178 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_489
timestamp 1607639953
transform 1 0 46074 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_498
timestamp 1607639953
transform 1 0 46902 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_486
timestamp 1607639953
transform 1 0 45798 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1607639953
transform 1 0 45982 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_525
timestamp 1607639953
transform 1 0 49386 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_513
timestamp 1607639953
transform 1 0 48282 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_520
timestamp 1607639953
transform 1 0 48926 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_518
timestamp 1607639953
transform 1 0 48742 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_510
timestamp 1607639953
transform 1 0 48006 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1607639953
transform 1 0 48834 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_550
timestamp 1607639953
transform 1 0 51686 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_537
timestamp 1607639953
transform 1 0 50490 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_544
timestamp 1607639953
transform 1 0 51134 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_532
timestamp 1607639953
transform 1 0 50030 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1607639953
transform 1 0 51594 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_562
timestamp 1607639953
transform 1 0 52790 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_568
timestamp 1607639953
transform 1 0 53342 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_556
timestamp 1607639953
transform 1 0 52238 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_586
timestamp 1607639953
transform 1 0 54998 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_574
timestamp 1607639953
transform 1 0 53894 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_593
timestamp 1607639953
transform 1 0 55642 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_581
timestamp 1607639953
transform 1 0 54538 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1607639953
transform 1 0 54446 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_611
timestamp 1607639953
transform 1 0 57298 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_598
timestamp 1607639953
transform 1 0 56102 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_605
timestamp 1607639953
transform 1 0 56746 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1607639953
transform 1 0 57206 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_623
timestamp 1607639953
transform 1 0 58402 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_617
timestamp 1607639953
transform 1 0 57850 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1607639953
transform -1 0 58862 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1607639953
transform -1 0 58862 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1607639953
transform 1 0 2466 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1607639953
transform 1 0 1362 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1607639953
transform 1 0 1086 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_44
timestamp 1607639953
transform 1 0 5134 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1607639953
transform 1 0 4030 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1607639953
transform 1 0 3570 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1607639953
transform 1 0 3938 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_60
timestamp 1607639953
transform 1 0 6606 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_48
timestamp 1607639953
transform 1 0 5502 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _122_
timestamp 1607639953
transform 1 0 5226 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_84
timestamp 1607639953
transform 1 0 8814 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_72
timestamp 1607639953
transform 1 0 7710 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1607639953
transform 1 0 10746 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1607639953
transform 1 0 9642 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1607639953
transform 1 0 9550 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1607639953
transform 1 0 12954 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1607639953
transform 1 0 11850 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1607639953
transform 1 0 15254 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1607639953
transform 1 0 14058 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1607639953
transform 1 0 15162 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1607639953
transform 1 0 16358 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1607639953
transform 1 0 18566 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1607639953
transform 1 0 17462 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1607639953
transform 1 0 20866 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1607639953
transform 1 0 19670 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1607639953
transform 1 0 20774 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1607639953
transform 1 0 23074 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1607639953
transform 1 0 21970 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1607639953
transform 1 0 25282 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1607639953
transform 1 0 24178 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_276
timestamp 1607639953
transform 1 0 26478 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1607639953
transform 1 0 26386 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_300
timestamp 1607639953
transform 1 0 28686 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_288
timestamp 1607639953
transform 1 0 27582 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_324
timestamp 1607639953
transform 1 0 30894 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_312
timestamp 1607639953
transform 1 0 29790 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_349
timestamp 1607639953
transform 1 0 33194 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_337
timestamp 1607639953
transform 1 0 32090 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1607639953
transform 1 0 31998 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_373
timestamp 1607639953
transform 1 0 35402 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_361
timestamp 1607639953
transform 1 0 34298 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_385
timestamp 1607639953
transform 1 0 36506 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_410
timestamp 1607639953
transform 1 0 38806 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_398
timestamp 1607639953
transform 1 0 37702 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1607639953
transform 1 0 37610 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_434
timestamp 1607639953
transform 1 0 41014 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_422
timestamp 1607639953
transform 1 0 39910 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_459
timestamp 1607639953
transform 1 0 43314 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_446
timestamp 1607639953
transform 1 0 42118 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1607639953
transform 1 0 43222 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_483
timestamp 1607639953
transform 1 0 45522 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_471
timestamp 1607639953
transform 1 0 44418 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_495
timestamp 1607639953
transform 1 0 46626 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_520
timestamp 1607639953
transform 1 0 48926 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_507
timestamp 1607639953
transform 1 0 47730 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1607639953
transform 1 0 48834 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_544
timestamp 1607639953
transform 1 0 51134 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_532
timestamp 1607639953
transform 1 0 50030 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_568
timestamp 1607639953
transform 1 0 53342 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_556
timestamp 1607639953
transform 1 0 52238 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_593
timestamp 1607639953
transform 1 0 55642 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_581
timestamp 1607639953
transform 1 0 54538 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1607639953
transform 1 0 54446 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_605
timestamp 1607639953
transform 1 0 56746 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_617
timestamp 1607639953
transform 1 0 57850 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1607639953
transform -1 0 58862 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1607639953
transform 1 0 2466 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1607639953
transform 1 0 1362 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1607639953
transform 1 0 1086 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1607639953
transform 1 0 4674 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1607639953
transform 1 0 3570 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1607639953
transform 1 0 6790 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1607639953
transform 1 0 6514 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1607639953
transform 1 0 5778 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1607639953
transform 1 0 6698 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_82
timestamp 1607639953
transform 1 0 8630 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_74
timestamp 1607639953
transform 1 0 7894 0 1 7072
box -38 -48 222 592
use BUFX2  BUFX2
timestamp 1608122862
transform 1 0 8078 0 1 7072
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_9_106
timestamp 1607639953
transform 1 0 10838 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_94
timestamp 1607639953
transform 1 0 9734 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1607639953
transform 1 0 12402 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1607639953
transform 1 0 11942 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1607639953
transform 1 0 12310 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_153
timestamp 1607639953
transform 1 0 15162 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_141
timestamp 1607639953
transform 1 0 14058 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_135
timestamp 1607639953
transform 1 0 13506 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _069_
timestamp 1607639953
transform 1 0 13782 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_165
timestamp 1607639953
transform 1 0 16266 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1607639953
transform 1 0 19118 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1607639953
transform 1 0 18014 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_177
timestamp 1607639953
transform 1 0 17370 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1607639953
transform 1 0 17922 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1607639953
transform 1 0 21326 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1607639953
transform 1 0 20222 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1607639953
transform 1 0 22430 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1607639953
transform 1 0 24730 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1607639953
transform 1 0 23626 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1607639953
transform 1 0 23534 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1607639953
transform 1 0 26938 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_269
timestamp 1607639953
transform 1 0 25834 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_306
timestamp 1607639953
transform 1 0 29238 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1607639953
transform 1 0 28042 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1607639953
transform 1 0 29146 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_330
timestamp 1607639953
transform 1 0 31446 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_318
timestamp 1607639953
transform 1 0 30342 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_342
timestamp 1607639953
transform 1 0 32550 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_367
timestamp 1607639953
transform 1 0 34850 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_354
timestamp 1607639953
transform 1 0 33654 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1607639953
transform 1 0 34758 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_391
timestamp 1607639953
transform 1 0 37058 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_379
timestamp 1607639953
transform 1 0 35954 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_415
timestamp 1607639953
transform 1 0 39266 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_403
timestamp 1607639953
transform 1 0 38162 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_440
timestamp 1607639953
transform 1 0 41566 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_428
timestamp 1607639953
transform 1 0 40462 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1607639953
transform 1 0 40370 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_452
timestamp 1607639953
transform 1 0 42670 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_476
timestamp 1607639953
transform 1 0 44878 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_464
timestamp 1607639953
transform 1 0 43774 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_501
timestamp 1607639953
transform 1 0 47178 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_489
timestamp 1607639953
transform 1 0 46074 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1607639953
transform 1 0 45982 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_525
timestamp 1607639953
transform 1 0 49386 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_513
timestamp 1607639953
transform 1 0 48282 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_550
timestamp 1607639953
transform 1 0 51686 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_537
timestamp 1607639953
transform 1 0 50490 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1607639953
transform 1 0 51594 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_562
timestamp 1607639953
transform 1 0 52790 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_586
timestamp 1607639953
transform 1 0 54998 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_574
timestamp 1607639953
transform 1 0 53894 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_611
timestamp 1607639953
transform 1 0 57298 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_598
timestamp 1607639953
transform 1 0 56102 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1607639953
transform 1 0 57206 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_623
timestamp 1607639953
transform 1 0 58402 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1607639953
transform -1 0 58862 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1607639953
transform 1 0 2466 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1607639953
transform 1 0 1362 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1607639953
transform 1 0 1086 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1607639953
transform 1 0 5134 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1607639953
transform 1 0 4030 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1607639953
transform 1 0 3570 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1607639953
transform 1 0 3938 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1607639953
transform 1 0 6238 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1607639953
transform 1 0 8446 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1607639953
transform 1 0 7342 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1607639953
transform 1 0 10746 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1607639953
transform 1 0 9642 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1607639953
transform 1 0 9550 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1607639953
transform 1 0 12954 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1607639953
transform 1 0 11850 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1607639953
transform 1 0 15254 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1607639953
transform 1 0 14058 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1607639953
transform 1 0 15162 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1607639953
transform 1 0 16358 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1607639953
transform 1 0 18566 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1607639953
transform 1 0 17462 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1607639953
transform 1 0 20866 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1607639953
transform 1 0 19670 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1607639953
transform 1 0 20774 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1607639953
transform 1 0 23074 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1607639953
transform 1 0 21970 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_262
timestamp 1607639953
transform 1 0 25190 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_251
timestamp 1607639953
transform 1 0 24178 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _104_
timestamp 1607639953
transform 1 0 24914 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_276
timestamp 1607639953
transform 1 0 26478 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_274
timestamp 1607639953
transform 1 0 26294 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1607639953
transform 1 0 26386 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_300
timestamp 1607639953
transform 1 0 28686 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_288
timestamp 1607639953
transform 1 0 27582 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_324
timestamp 1607639953
transform 1 0 30894 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_312
timestamp 1607639953
transform 1 0 29790 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_349
timestamp 1607639953
transform 1 0 33194 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_337
timestamp 1607639953
transform 1 0 32090 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1607639953
transform 1 0 31998 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_373
timestamp 1607639953
transform 1 0 35402 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_361
timestamp 1607639953
transform 1 0 34298 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_385
timestamp 1607639953
transform 1 0 36506 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_410
timestamp 1607639953
transform 1 0 38806 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_398
timestamp 1607639953
transform 1 0 37702 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1607639953
transform 1 0 37610 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_434
timestamp 1607639953
transform 1 0 41014 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_422
timestamp 1607639953
transform 1 0 39910 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_459
timestamp 1607639953
transform 1 0 43314 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_446
timestamp 1607639953
transform 1 0 42118 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1607639953
transform 1 0 43222 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_483
timestamp 1607639953
transform 1 0 45522 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_471
timestamp 1607639953
transform 1 0 44418 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_504
timestamp 1607639953
transform 1 0 47454 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_492
timestamp 1607639953
transform 1 0 46350 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _094_
timestamp 1607639953
transform 1 0 46074 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_525
timestamp 1607639953
transform 1 0 49386 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_520
timestamp 1607639953
transform 1 0 48926 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_516
timestamp 1607639953
transform 1 0 48558 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1607639953
transform 1 0 48834 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1607639953
transform 1 0 49110 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_549
timestamp 1607639953
transform 1 0 51594 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_537
timestamp 1607639953
transform 1 0 50490 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_561
timestamp 1607639953
transform 1 0 52698 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_593
timestamp 1607639953
transform 1 0 55642 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_581
timestamp 1607639953
transform 1 0 54538 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_579
timestamp 1607639953
transform 1 0 54354 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_573
timestamp 1607639953
transform 1 0 53802 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1607639953
transform 1 0 54446 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_605
timestamp 1607639953
transform 1 0 56746 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_617
timestamp 1607639953
transform 1 0 57850 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1607639953
transform -1 0 58862 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1607639953
transform 1 0 2466 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1607639953
transform 1 0 1362 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1607639953
transform 1 0 1086 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_34
timestamp 1607639953
transform 1 0 4214 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1607639953
transform 1 0 3570 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _021_
timestamp 1607639953
transform 1 0 3938 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1607639953
transform 1 0 6790 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_58
timestamp 1607639953
transform 1 0 6422 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_46
timestamp 1607639953
transform 1 0 5318 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1607639953
transform 1 0 6698 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_84
timestamp 1607639953
transform 1 0 8814 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_74
timestamp 1607639953
transform 1 0 7894 0 1 8160
box -38 -48 222 592
use BUFX4  BUFX4
timestamp 1608122862
transform 1 0 8078 0 1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_11_108
timestamp 1607639953
transform 1 0 11022 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_96
timestamp 1607639953
transform 1 0 9918 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1607639953
transform 1 0 12402 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1607639953
transform 1 0 12126 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1607639953
transform 1 0 12310 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1607639953
transform 1 0 14610 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1607639953
transform 1 0 13506 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1607639953
transform 1 0 16818 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1607639953
transform 1 0 15714 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1607639953
transform 1 0 19118 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1607639953
transform 1 0 18014 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1607639953
transform 1 0 17922 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1607639953
transform 1 0 21326 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1607639953
transform 1 0 20222 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1607639953
transform 1 0 22430 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1607639953
transform 1 0 24730 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1607639953
transform 1 0 23626 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1607639953
transform 1 0 23534 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1607639953
transform 1 0 26938 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_269
timestamp 1607639953
transform 1 0 25834 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_306
timestamp 1607639953
transform 1 0 29238 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1607639953
transform 1 0 28042 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1607639953
transform 1 0 29146 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_330
timestamp 1607639953
transform 1 0 31446 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_318
timestamp 1607639953
transform 1 0 30342 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_342
timestamp 1607639953
transform 1 0 32550 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_367
timestamp 1607639953
transform 1 0 34850 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_354
timestamp 1607639953
transform 1 0 33654 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1607639953
transform 1 0 34758 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_391
timestamp 1607639953
transform 1 0 37058 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_379
timestamp 1607639953
transform 1 0 35954 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_415
timestamp 1607639953
transform 1 0 39266 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_403
timestamp 1607639953
transform 1 0 38162 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_440
timestamp 1607639953
transform 1 0 41566 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_428
timestamp 1607639953
transform 1 0 40462 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_426
timestamp 1607639953
transform 1 0 40278 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_422
timestamp 1607639953
transform 1 0 39910 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1607639953
transform 1 0 40370 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _080_
timestamp 1607639953
transform 1 0 39634 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_452
timestamp 1607639953
transform 1 0 42670 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_476
timestamp 1607639953
transform 1 0 44878 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_464
timestamp 1607639953
transform 1 0 43774 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_501
timestamp 1607639953
transform 1 0 47178 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_497
timestamp 1607639953
transform 1 0 46810 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_489
timestamp 1607639953
transform 1 0 46074 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1607639953
transform 1 0 45982 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _200_
timestamp 1607639953
transform 1 0 46902 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_527
timestamp 1607639953
transform 1 0 49570 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_515
timestamp 1607639953
transform 1 0 48466 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_509
timestamp 1607639953
transform 1 0 47914 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _178_
timestamp 1607639953
transform 1 0 48190 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_550
timestamp 1607639953
transform 1 0 51686 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_547
timestamp 1607639953
transform 1 0 51410 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_539
timestamp 1607639953
transform 1 0 50674 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1607639953
transform 1 0 51594 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_562
timestamp 1607639953
transform 1 0 52790 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_586
timestamp 1607639953
transform 1 0 54998 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_574
timestamp 1607639953
transform 1 0 53894 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_611
timestamp 1607639953
transform 1 0 57298 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_598
timestamp 1607639953
transform 1 0 56102 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1607639953
transform 1 0 57206 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_623
timestamp 1607639953
transform 1 0 58402 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1607639953
transform -1 0 58862 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1607639953
transform 1 0 2466 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1607639953
transform 1 0 1362 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1607639953
transform 1 0 1086 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1607639953
transform 1 0 5134 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1607639953
transform 1 0 4030 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1607639953
transform 1 0 3570 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1607639953
transform 1 0 3938 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1607639953
transform 1 0 6238 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1607639953
transform 1 0 8446 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1607639953
transform 1 0 7342 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1607639953
transform 1 0 10746 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1607639953
transform 1 0 9642 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1607639953
transform 1 0 9550 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1607639953
transform 1 0 12954 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1607639953
transform 1 0 11850 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1607639953
transform 1 0 15254 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1607639953
transform 1 0 14058 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1607639953
transform 1 0 15162 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1607639953
transform 1 0 16358 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1607639953
transform 1 0 18566 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1607639953
transform 1 0 17462 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1607639953
transform 1 0 20866 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1607639953
transform 1 0 19670 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1607639953
transform 1 0 20774 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1607639953
transform 1 0 23074 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1607639953
transform 1 0 21970 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1607639953
transform 1 0 25282 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1607639953
transform 1 0 24178 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_276
timestamp 1607639953
transform 1 0 26478 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1607639953
transform 1 0 26386 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_300
timestamp 1607639953
transform 1 0 28686 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_288
timestamp 1607639953
transform 1 0 27582 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_324
timestamp 1607639953
transform 1 0 30894 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_312
timestamp 1607639953
transform 1 0 29790 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_349
timestamp 1607639953
transform 1 0 33194 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_337
timestamp 1607639953
transform 1 0 32090 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1607639953
transform 1 0 31998 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_373
timestamp 1607639953
transform 1 0 35402 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_361
timestamp 1607639953
transform 1 0 34298 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_385
timestamp 1607639953
transform 1 0 36506 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_410
timestamp 1607639953
transform 1 0 38806 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_398
timestamp 1607639953
transform 1 0 37702 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1607639953
transform 1 0 37610 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_434
timestamp 1607639953
transform 1 0 41014 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_422
timestamp 1607639953
transform 1 0 39910 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_459
timestamp 1607639953
transform 1 0 43314 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_446
timestamp 1607639953
transform 1 0 42118 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1607639953
transform 1 0 43222 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_483
timestamp 1607639953
transform 1 0 45522 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_471
timestamp 1607639953
transform 1 0 44418 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_495
timestamp 1607639953
transform 1 0 46626 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_520
timestamp 1607639953
transform 1 0 48926 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_507
timestamp 1607639953
transform 1 0 47730 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1607639953
transform 1 0 48834 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_544
timestamp 1607639953
transform 1 0 51134 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_532
timestamp 1607639953
transform 1 0 50030 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_568
timestamp 1607639953
transform 1 0 53342 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_556
timestamp 1607639953
transform 1 0 52238 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_593
timestamp 1607639953
transform 1 0 55642 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_581
timestamp 1607639953
transform 1 0 54538 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1607639953
transform 1 0 54446 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_605
timestamp 1607639953
transform 1 0 56746 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_617
timestamp 1607639953
transform 1 0 57850 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1607639953
transform -1 0 58862 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1607639953
transform 1 0 2466 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1607639953
transform 1 0 1362 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1607639953
transform 1 0 2466 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1607639953
transform 1 0 1362 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1607639953
transform 1 0 1086 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1607639953
transform 1 0 1086 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1607639953
transform 1 0 5134 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1607639953
transform 1 0 4030 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1607639953
transform 1 0 3570 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1607639953
transform 1 0 4674 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1607639953
transform 1 0 3570 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1607639953
transform 1 0 3938 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1607639953
transform 1 0 6238 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1607639953
transform 1 0 6790 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1607639953
transform 1 0 6514 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1607639953
transform 1 0 5778 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1607639953
transform 1 0 6698 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1607639953
transform 1 0 8446 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1607639953
transform 1 0 7342 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_74
timestamp 1607639953
transform 1 0 7894 0 1 9248
box -38 -48 222 592
use CLKBUF1  CLKBUF1
timestamp 1608122862
transform 1 0 8078 0 1 9248
box 0 -48 1656 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1607639953
transform 1 0 10746 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1607639953
transform 1 0 9642 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_110
timestamp 1607639953
transform 1 0 11206 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1607639953
transform 1 0 10102 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_94
timestamp 1607639953
transform 1 0 9734 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1607639953
transform 1 0 9550 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _125_
timestamp 1607639953
transform 1 0 9826 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_129
timestamp 1607639953
transform 1 0 12954 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1607639953
transform 1 0 11850 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1607639953
transform 1 0 12402 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1607639953
transform 1 0 12310 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1607639953
transform 1 0 15254 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1607639953
transform 1 0 14058 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1607639953
transform 1 0 14610 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1607639953
transform 1 0 13506 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1607639953
transform 1 0 15162 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1607639953
transform 1 0 16358 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1607639953
transform 1 0 16818 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1607639953
transform 1 0 15714 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1607639953
transform 1 0 18566 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1607639953
transform 1 0 17462 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1607639953
transform 1 0 19118 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1607639953
transform 1 0 18014 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1607639953
transform 1 0 17922 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1607639953
transform 1 0 20866 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1607639953
transform 1 0 19670 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_215
timestamp 1607639953
transform 1 0 20866 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_208
timestamp 1607639953
transform 1 0 20222 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1607639953
transform 1 0 20774 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _190_
timestamp 1607639953
transform 1 0 20590 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1607639953
transform 1 0 23074 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1607639953
transform 1 0 21970 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_239
timestamp 1607639953
transform 1 0 23074 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_227
timestamp 1607639953
transform 1 0 21970 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1607639953
transform 1 0 25282 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1607639953
transform 1 0 24178 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1607639953
transform 1 0 24730 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1607639953
transform 1 0 23626 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 1607639953
transform 1 0 23442 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1607639953
transform 1 0 23534 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_276
timestamp 1607639953
transform 1 0 26478 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1607639953
transform 1 0 26938 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_269
timestamp 1607639953
transform 1 0 25834 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1607639953
transform 1 0 26386 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_300
timestamp 1607639953
transform 1 0 28686 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_288
timestamp 1607639953
transform 1 0 27582 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_306
timestamp 1607639953
transform 1 0 29238 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1607639953
transform 1 0 28042 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1607639953
transform 1 0 29146 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_324
timestamp 1607639953
transform 1 0 30894 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_312
timestamp 1607639953
transform 1 0 29790 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_330
timestamp 1607639953
transform 1 0 31446 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_318
timestamp 1607639953
transform 1 0 30342 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_345
timestamp 1607639953
transform 1 0 32826 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_340
timestamp 1607639953
transform 1 0 32366 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_342
timestamp 1607639953
transform 1 0 32550 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1607639953
transform 1 0 31998 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1607639953
transform 1 0 32090 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _015_
timestamp 1607639953
transform 1 0 32550 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_368
timestamp 1607639953
transform 1 0 34942 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_356
timestamp 1607639953
transform 1 0 33838 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_367
timestamp 1607639953
transform 1 0 34850 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_354
timestamp 1607639953
transform 1 0 33654 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1607639953
transform 1 0 34758 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1607639953
transform 1 0 33562 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_396
timestamp 1607639953
transform 1 0 37518 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_392
timestamp 1607639953
transform 1 0 37150 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_380
timestamp 1607639953
transform 1 0 36046 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_391
timestamp 1607639953
transform 1 0 37058 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_379
timestamp 1607639953
transform 1 0 35954 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_410
timestamp 1607639953
transform 1 0 38806 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_398
timestamp 1607639953
transform 1 0 37702 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_415
timestamp 1607639953
transform 1 0 39266 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_403
timestamp 1607639953
transform 1 0 38162 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1607639953
transform 1 0 37610 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_434
timestamp 1607639953
transform 1 0 41014 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_422
timestamp 1607639953
transform 1 0 39910 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_440
timestamp 1607639953
transform 1 0 41566 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_428
timestamp 1607639953
transform 1 0 40462 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1607639953
transform 1 0 40370 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_459
timestamp 1607639953
transform 1 0 43314 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_446
timestamp 1607639953
transform 1 0 42118 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_452
timestamp 1607639953
transform 1 0 42670 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1607639953
transform 1 0 43222 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_483
timestamp 1607639953
transform 1 0 45522 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_471
timestamp 1607639953
transform 1 0 44418 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_476
timestamp 1607639953
transform 1 0 44878 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_464
timestamp 1607639953
transform 1 0 43774 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_495
timestamp 1607639953
transform 1 0 46626 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_501
timestamp 1607639953
transform 1 0 47178 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_489
timestamp 1607639953
transform 1 0 46074 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1607639953
transform 1 0 45982 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_523
timestamp 1607639953
transform 1 0 49202 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_507
timestamp 1607639953
transform 1 0 47730 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_525
timestamp 1607639953
transform 1 0 49386 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_513
timestamp 1607639953
transform 1 0 48282 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1607639953
transform 1 0 48834 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _159_
timestamp 1607639953
transform 1 0 48926 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_547
timestamp 1607639953
transform 1 0 51410 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_535
timestamp 1607639953
transform 1 0 50306 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_550
timestamp 1607639953
transform 1 0 51686 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_537
timestamp 1607639953
transform 1 0 50490 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1607639953
transform 1 0 51594 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_571
timestamp 1607639953
transform 1 0 53618 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_559
timestamp 1607639953
transform 1 0 52514 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_562
timestamp 1607639953
transform 1 0 52790 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_593
timestamp 1607639953
transform 1 0 55642 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_581
timestamp 1607639953
transform 1 0 54538 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_579
timestamp 1607639953
transform 1 0 54354 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_586
timestamp 1607639953
transform 1 0 54998 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_574
timestamp 1607639953
transform 1 0 53894 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1607639953
transform 1 0 54446 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_605
timestamp 1607639953
transform 1 0 56746 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_611
timestamp 1607639953
transform 1 0 57298 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_598
timestamp 1607639953
transform 1 0 56102 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1607639953
transform 1 0 57206 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_617
timestamp 1607639953
transform 1 0 57850 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_623
timestamp 1607639953
transform 1 0 58402 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1607639953
transform -1 0 58862 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1607639953
transform -1 0 58862 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1607639953
transform 1 0 2466 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1607639953
transform 1 0 1362 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1607639953
transform 1 0 1086 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1607639953
transform 1 0 4674 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1607639953
transform 1 0 3570 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1607639953
transform 1 0 6790 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1607639953
transform 1 0 6514 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1607639953
transform 1 0 5778 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1607639953
transform 1 0 6698 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_74
timestamp 1607639953
transform 1 0 7894 0 1 10336
box -38 -48 222 592
use HAX1  HAX1
timestamp 1608122862
transform 1 0 8078 0 1 10336
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1607639953
transform 1 0 11206 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1607639953
transform 1 0 10102 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1607639953
transform 1 0 12402 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1607639953
transform 1 0 12310 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1607639953
transform 1 0 14610 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1607639953
transform 1 0 13506 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_171
timestamp 1607639953
transform 1 0 16818 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_159
timestamp 1607639953
transform 1 0 15714 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1607639953
transform 1 0 19118 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1607639953
transform 1 0 18014 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1607639953
transform 1 0 17922 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_220
timestamp 1607639953
transform 1 0 21326 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1607639953
transform 1 0 20222 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_232
timestamp 1607639953
transform 1 0 22430 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1607639953
transform 1 0 24730 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1607639953
transform 1 0 23626 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1607639953
transform 1 0 23534 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1607639953
transform 1 0 26938 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_269
timestamp 1607639953
transform 1 0 25834 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_306
timestamp 1607639953
transform 1 0 29238 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1607639953
transform 1 0 28042 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1607639953
transform 1 0 29146 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_325
timestamp 1607639953
transform 1 0 30986 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_313
timestamp 1607639953
transform 1 0 29882 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1607639953
transform 1 0 29606 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1607639953
transform 1 0 33194 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1607639953
transform 1 0 32090 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_367
timestamp 1607639953
transform 1 0 34850 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_365
timestamp 1607639953
transform 1 0 34666 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_361
timestamp 1607639953
transform 1 0 34298 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1607639953
transform 1 0 34758 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_391
timestamp 1607639953
transform 1 0 37058 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_379
timestamp 1607639953
transform 1 0 35954 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_415
timestamp 1607639953
transform 1 0 39266 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_403
timestamp 1607639953
transform 1 0 38162 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_440
timestamp 1607639953
transform 1 0 41566 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_428
timestamp 1607639953
transform 1 0 40462 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1607639953
transform 1 0 40370 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_452
timestamp 1607639953
transform 1 0 42670 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_476
timestamp 1607639953
transform 1 0 44878 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_464
timestamp 1607639953
transform 1 0 43774 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_501
timestamp 1607639953
transform 1 0 47178 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_489
timestamp 1607639953
transform 1 0 46074 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1607639953
transform 1 0 45982 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_525
timestamp 1607639953
transform 1 0 49386 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_513
timestamp 1607639953
transform 1 0 48282 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_550
timestamp 1607639953
transform 1 0 51686 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_537
timestamp 1607639953
transform 1 0 50490 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1607639953
transform 1 0 51594 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_562
timestamp 1607639953
transform 1 0 52790 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_586
timestamp 1607639953
transform 1 0 54998 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_574
timestamp 1607639953
transform 1 0 53894 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_611
timestamp 1607639953
transform 1 0 57298 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_598
timestamp 1607639953
transform 1 0 56102 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1607639953
transform 1 0 57206 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_623
timestamp 1607639953
transform 1 0 58402 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1607639953
transform -1 0 58862 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1607639953
transform 1 0 2466 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1607639953
transform 1 0 1362 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1607639953
transform 1 0 1086 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1607639953
transform 1 0 5134 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1607639953
transform 1 0 4030 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1607639953
transform 1 0 3570 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1607639953
transform 1 0 3938 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1607639953
transform 1 0 6238 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1607639953
transform 1 0 8446 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1607639953
transform 1 0 7342 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1607639953
transform 1 0 10746 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1607639953
transform 1 0 9642 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1607639953
transform 1 0 9550 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_129
timestamp 1607639953
transform 1 0 12954 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1607639953
transform 1 0 11850 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1607639953
transform 1 0 15254 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1607639953
transform 1 0 14058 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1607639953
transform 1 0 15162 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1607639953
transform 1 0 16358 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_190
timestamp 1607639953
transform 1 0 18566 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1607639953
transform 1 0 17462 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1607639953
transform 1 0 20866 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1607639953
transform 1 0 19670 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1607639953
transform 1 0 20774 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1607639953
transform 1 0 23074 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1607639953
transform 1 0 21970 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1607639953
transform 1 0 25282 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1607639953
transform 1 0 24178 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_276
timestamp 1607639953
transform 1 0 26478 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1607639953
transform 1 0 26386 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_300
timestamp 1607639953
transform 1 0 28686 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_288
timestamp 1607639953
transform 1 0 27582 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_324
timestamp 1607639953
transform 1 0 30894 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_312
timestamp 1607639953
transform 1 0 29790 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_349
timestamp 1607639953
transform 1 0 33194 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_337
timestamp 1607639953
transform 1 0 32090 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1607639953
transform 1 0 31998 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_373
timestamp 1607639953
transform 1 0 35402 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_361
timestamp 1607639953
transform 1 0 34298 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_385
timestamp 1607639953
transform 1 0 36506 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_410
timestamp 1607639953
transform 1 0 38806 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_398
timestamp 1607639953
transform 1 0 37702 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1607639953
transform 1 0 37610 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_434
timestamp 1607639953
transform 1 0 41014 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_422
timestamp 1607639953
transform 1 0 39910 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_459
timestamp 1607639953
transform 1 0 43314 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_446
timestamp 1607639953
transform 1 0 42118 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1607639953
transform 1 0 43222 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_483
timestamp 1607639953
transform 1 0 45522 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_471
timestamp 1607639953
transform 1 0 44418 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_495
timestamp 1607639953
transform 1 0 46626 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_520
timestamp 1607639953
transform 1 0 48926 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_507
timestamp 1607639953
transform 1 0 47730 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1607639953
transform 1 0 48834 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_544
timestamp 1607639953
transform 1 0 51134 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_532
timestamp 1607639953
transform 1 0 50030 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_568
timestamp 1607639953
transform 1 0 53342 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_556
timestamp 1607639953
transform 1 0 52238 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_593
timestamp 1607639953
transform 1 0 55642 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_581
timestamp 1607639953
transform 1 0 54538 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1607639953
transform 1 0 54446 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_605
timestamp 1607639953
transform 1 0 56746 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_617
timestamp 1607639953
transform 1 0 57850 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1607639953
transform -1 0 58862 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1607639953
transform 1 0 2466 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1607639953
transform 1 0 1362 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1607639953
transform 1 0 1086 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1607639953
transform 1 0 4674 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1607639953
transform 1 0 3570 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1607639953
transform 1 0 6790 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1607639953
transform 1 0 6514 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1607639953
transform 1 0 5778 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1607639953
transform 1 0 6698 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_80
timestamp 1607639953
transform 1 0 8446 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_74
timestamp 1607639953
transform 1 0 7894 0 1 11424
box -38 -48 222 592
use INV  INV
timestamp 1608122862
transform 1 0 8078 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_17_104
timestamp 1607639953
transform 1 0 10654 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_92
timestamp 1607639953
transform 1 0 9550 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1607639953
transform 1 0 12402 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_116
timestamp 1607639953
transform 1 0 11758 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1607639953
transform 1 0 12310 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1607639953
transform 1 0 14610 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1607639953
transform 1 0 13506 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_171
timestamp 1607639953
transform 1 0 16818 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_159
timestamp 1607639953
transform 1 0 15714 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1607639953
transform 1 0 19118 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_192
timestamp 1607639953
transform 1 0 18750 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_184
timestamp 1607639953
transform 1 0 18014 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1607639953
transform 1 0 17922 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _194_
timestamp 1607639953
transform 1 0 18842 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_220
timestamp 1607639953
transform 1 0 21326 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1607639953
transform 1 0 20222 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_232
timestamp 1607639953
transform 1 0 22430 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1607639953
transform 1 0 24730 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1607639953
transform 1 0 23626 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1607639953
transform 1 0 23534 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1607639953
transform 1 0 26938 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_269
timestamp 1607639953
transform 1 0 25834 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_306
timestamp 1607639953
transform 1 0 29238 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1607639953
transform 1 0 28042 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1607639953
transform 1 0 29146 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_330
timestamp 1607639953
transform 1 0 31446 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_318
timestamp 1607639953
transform 1 0 30342 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_342
timestamp 1607639953
transform 1 0 32550 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_367
timestamp 1607639953
transform 1 0 34850 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_354
timestamp 1607639953
transform 1 0 33654 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1607639953
transform 1 0 34758 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_391
timestamp 1607639953
transform 1 0 37058 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_379
timestamp 1607639953
transform 1 0 35954 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_415
timestamp 1607639953
transform 1 0 39266 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_403
timestamp 1607639953
transform 1 0 38162 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_440
timestamp 1607639953
transform 1 0 41566 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_428
timestamp 1607639953
transform 1 0 40462 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1607639953
transform 1 0 40370 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_452
timestamp 1607639953
transform 1 0 42670 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_476
timestamp 1607639953
transform 1 0 44878 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_464
timestamp 1607639953
transform 1 0 43774 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_501
timestamp 1607639953
transform 1 0 47178 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_489
timestamp 1607639953
transform 1 0 46074 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1607639953
transform 1 0 45982 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_526
timestamp 1607639953
transform 1 0 49478 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_521
timestamp 1607639953
transform 1 0 49018 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_513
timestamp 1607639953
transform 1 0 48282 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _169_
timestamp 1607639953
transform 1 0 49202 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_550
timestamp 1607639953
transform 1 0 51686 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_546
timestamp 1607639953
transform 1 0 51318 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_538
timestamp 1607639953
transform 1 0 50582 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1607639953
transform 1 0 51594 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_562
timestamp 1607639953
transform 1 0 52790 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_586
timestamp 1607639953
transform 1 0 54998 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_574
timestamp 1607639953
transform 1 0 53894 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _172_
timestamp 1607639953
transform 1 0 55734 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_611
timestamp 1607639953
transform 1 0 57298 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_609
timestamp 1607639953
transform 1 0 57114 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_597
timestamp 1607639953
transform 1 0 56010 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1607639953
transform 1 0 57206 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_623
timestamp 1607639953
transform 1 0 58402 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1607639953
transform -1 0 58862 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1607639953
transform 1 0 2466 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1607639953
transform 1 0 1362 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1607639953
transform 1 0 1086 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1607639953
transform 1 0 5134 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1607639953
transform 1 0 4030 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1607639953
transform 1 0 3570 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1607639953
transform 1 0 3938 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1607639953
transform 1 0 6238 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1607639953
transform 1 0 8446 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1607639953
transform 1 0 7342 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1607639953
transform 1 0 10746 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1607639953
transform 1 0 9642 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1607639953
transform 1 0 9550 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1607639953
transform 1 0 12954 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1607639953
transform 1 0 11850 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1607639953
transform 1 0 15254 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1607639953
transform 1 0 14058 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1607639953
transform 1 0 15162 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1607639953
transform 1 0 16358 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1607639953
transform 1 0 18566 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1607639953
transform 1 0 17462 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1607639953
transform 1 0 20866 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1607639953
transform 1 0 20590 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_208
timestamp 1607639953
transform 1 0 20222 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_202
timestamp 1607639953
transform 1 0 19670 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1607639953
transform 1 0 20774 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _001_
timestamp 1607639953
transform 1 0 20314 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1607639953
transform 1 0 23074 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1607639953
transform 1 0 21970 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_256
timestamp 1607639953
transform 1 0 24638 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_251
timestamp 1607639953
transform 1 0 24178 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _017_
timestamp 1607639953
transform 1 0 24362 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_276
timestamp 1607639953
transform 1 0 26478 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_274
timestamp 1607639953
transform 1 0 26294 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_268
timestamp 1607639953
transform 1 0 25742 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1607639953
transform 1 0 26386 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_300
timestamp 1607639953
transform 1 0 28686 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_288
timestamp 1607639953
transform 1 0 27582 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_324
timestamp 1607639953
transform 1 0 30894 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_312
timestamp 1607639953
transform 1 0 29790 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_351
timestamp 1607639953
transform 1 0 33378 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_345
timestamp 1607639953
transform 1 0 32826 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_337
timestamp 1607639953
transform 1 0 32090 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1607639953
transform 1 0 31998 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _154_
timestamp 1607639953
transform 1 0 33102 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_363
timestamp 1607639953
transform 1 0 34482 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_395
timestamp 1607639953
transform 1 0 37426 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_387
timestamp 1607639953
transform 1 0 36690 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_375
timestamp 1607639953
transform 1 0 35586 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_410
timestamp 1607639953
transform 1 0 38806 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_398
timestamp 1607639953
transform 1 0 37702 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1607639953
transform 1 0 37610 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_434
timestamp 1607639953
transform 1 0 41014 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_422
timestamp 1607639953
transform 1 0 39910 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_459
timestamp 1607639953
transform 1 0 43314 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_456
timestamp 1607639953
transform 1 0 43038 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_448
timestamp 1607639953
transform 1 0 42302 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_442
timestamp 1607639953
transform 1 0 41750 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1607639953
transform 1 0 43222 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _186_
timestamp 1607639953
transform 1 0 42026 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_484
timestamp 1607639953
transform 1 0 45614 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_472
timestamp 1607639953
transform 1 0 44510 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_467
timestamp 1607639953
transform 1 0 44050 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _129_
timestamp 1607639953
transform 1 0 44234 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_496
timestamp 1607639953
transform 1 0 46718 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_520
timestamp 1607639953
transform 1 0 48926 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_516
timestamp 1607639953
transform 1 0 48558 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_508
timestamp 1607639953
transform 1 0 47822 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1607639953
transform 1 0 48834 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_544
timestamp 1607639953
transform 1 0 51134 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_532
timestamp 1607639953
transform 1 0 50030 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_568
timestamp 1607639953
transform 1 0 53342 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_556
timestamp 1607639953
transform 1 0 52238 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_593
timestamp 1607639953
transform 1 0 55642 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_581
timestamp 1607639953
transform 1 0 54538 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1607639953
transform 1 0 54446 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_605
timestamp 1607639953
transform 1 0 56746 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_617
timestamp 1607639953
transform 1 0 57850 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1607639953
transform -1 0 58862 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1607639953
transform 1 0 2466 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1607639953
transform 1 0 1362 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1607639953
transform 1 0 2466 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1607639953
transform 1 0 1362 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1607639953
transform 1 0 1086 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1607639953
transform 1 0 1086 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1607639953
transform 1 0 5134 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1607639953
transform 1 0 4030 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1607639953
transform 1 0 3570 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1607639953
transform 1 0 4674 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1607639953
transform 1 0 3570 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1607639953
transform 1 0 3938 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1607639953
transform 1 0 6238 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1607639953
transform 1 0 6790 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1607639953
transform 1 0 6514 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1607639953
transform 1 0 5778 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1607639953
transform 1 0 6698 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1607639953
transform 1 0 8446 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1607639953
transform 1 0 7342 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_80
timestamp 1607639953
transform 1 0 8446 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_74
timestamp 1607639953
transform 1 0 7894 0 1 12512
box -38 -48 222 592
use INVX1  INVX1
timestamp 1608122862
transform 1 0 8078 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1607639953
transform 1 0 10746 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1607639953
transform 1 0 9642 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_104
timestamp 1607639953
transform 1 0 10654 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_92
timestamp 1607639953
transform 1 0 9550 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1607639953
transform 1 0 9550 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1607639953
transform 1 0 12954 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1607639953
transform 1 0 11850 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1607639953
transform 1 0 12402 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_116
timestamp 1607639953
transform 1 0 11758 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1607639953
transform 1 0 12310 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1607639953
transform 1 0 15254 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1607639953
transform 1 0 14058 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1607639953
transform 1 0 14610 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1607639953
transform 1 0 13506 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1607639953
transform 1 0 15162 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1607639953
transform 1 0 16358 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1607639953
transform 1 0 16818 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1607639953
transform 1 0 15714 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1607639953
transform 1 0 18566 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1607639953
transform 1 0 17462 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1607639953
transform 1 0 19118 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1607639953
transform 1 0 18014 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1607639953
transform 1 0 17922 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1607639953
transform 1 0 20866 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1607639953
transform 1 0 19670 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_220
timestamp 1607639953
transform 1 0 21326 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1607639953
transform 1 0 20222 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1607639953
transform 1 0 20774 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_239
timestamp 1607639953
transform 1 0 23074 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_227
timestamp 1607639953
transform 1 0 21970 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_242
timestamp 1607639953
transform 1 0 23350 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_230
timestamp 1607639953
transform 1 0 22246 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_226
timestamp 1607639953
transform 1 0 21878 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _197_
timestamp 1607639953
transform 1 0 21970 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_263
timestamp 1607639953
transform 1 0 25282 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_251
timestamp 1607639953
transform 1 0 24178 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_260
timestamp 1607639953
transform 1 0 25006 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_248
timestamp 1607639953
transform 1 0 23902 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1607639953
transform 1 0 23534 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _127_
timestamp 1607639953
transform 1 0 23626 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_276
timestamp 1607639953
transform 1 0 26478 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_284
timestamp 1607639953
transform 1 0 27214 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_272
timestamp 1607639953
transform 1 0 26110 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1607639953
transform 1 0 26386 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_300
timestamp 1607639953
transform 1 0 28686 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_288
timestamp 1607639953
transform 1 0 27582 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_306
timestamp 1607639953
transform 1 0 29238 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_303
timestamp 1607639953
transform 1 0 28962 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_291
timestamp 1607639953
transform 1 0 27858 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1607639953
transform 1 0 29146 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _181_
timestamp 1607639953
transform 1 0 27582 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_324
timestamp 1607639953
transform 1 0 30894 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_312
timestamp 1607639953
transform 1 0 29790 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_330
timestamp 1607639953
transform 1 0 31446 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_318
timestamp 1607639953
transform 1 0 30342 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_349
timestamp 1607639953
transform 1 0 33194 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_337
timestamp 1607639953
transform 1 0 32090 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_342
timestamp 1607639953
transform 1 0 32550 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1607639953
transform 1 0 31998 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_373
timestamp 1607639953
transform 1 0 35402 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_361
timestamp 1607639953
transform 1 0 34298 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_367
timestamp 1607639953
transform 1 0 34850 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_354
timestamp 1607639953
transform 1 0 33654 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1607639953
transform 1 0 34758 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_385
timestamp 1607639953
transform 1 0 36506 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_391
timestamp 1607639953
transform 1 0 37058 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_379
timestamp 1607639953
transform 1 0 35954 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_410
timestamp 1607639953
transform 1 0 38806 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_398
timestamp 1607639953
transform 1 0 37702 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_415
timestamp 1607639953
transform 1 0 39266 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_403
timestamp 1607639953
transform 1 0 38162 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1607639953
transform 1 0 37610 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_434
timestamp 1607639953
transform 1 0 41014 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_422
timestamp 1607639953
transform 1 0 39910 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_440
timestamp 1607639953
transform 1 0 41566 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_428
timestamp 1607639953
transform 1 0 40462 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1607639953
transform 1 0 40370 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_459
timestamp 1607639953
transform 1 0 43314 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_446
timestamp 1607639953
transform 1 0 42118 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_452
timestamp 1607639953
transform 1 0 42670 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1607639953
transform 1 0 43222 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_483
timestamp 1607639953
transform 1 0 45522 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_471
timestamp 1607639953
transform 1 0 44418 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_483
timestamp 1607639953
transform 1 0 45522 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_475
timestamp 1607639953
transform 1 0 44786 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_464
timestamp 1607639953
transform 1 0 43774 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _157_
timestamp 1607639953
transform 1 0 45614 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1607639953
transform 1 0 44510 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_495
timestamp 1607639953
transform 1 0 46626 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_501
timestamp 1607639953
transform 1 0 47178 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_489
timestamp 1607639953
transform 1 0 46074 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_487
timestamp 1607639953
transform 1 0 45890 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1607639953
transform 1 0 45982 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_520
timestamp 1607639953
transform 1 0 48926 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_507
timestamp 1607639953
transform 1 0 47730 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_525
timestamp 1607639953
transform 1 0 49386 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_513
timestamp 1607639953
transform 1 0 48282 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1607639953
transform 1 0 48834 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_544
timestamp 1607639953
transform 1 0 51134 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_532
timestamp 1607639953
transform 1 0 50030 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_550
timestamp 1607639953
transform 1 0 51686 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_537
timestamp 1607639953
transform 1 0 50490 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1607639953
transform 1 0 51594 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_568
timestamp 1607639953
transform 1 0 53342 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_556
timestamp 1607639953
transform 1 0 52238 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_564
timestamp 1607639953
transform 1 0 52974 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_558
timestamp 1607639953
transform 1 0 52422 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _075_
timestamp 1607639953
transform 1 0 52698 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_593
timestamp 1607639953
transform 1 0 55642 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_581
timestamp 1607639953
transform 1 0 54538 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_588
timestamp 1607639953
transform 1 0 55182 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_576
timestamp 1607639953
transform 1 0 54078 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1607639953
transform 1 0 54446 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_605
timestamp 1607639953
transform 1 0 56746 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_611
timestamp 1607639953
transform 1 0 57298 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_608
timestamp 1607639953
transform 1 0 57022 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_600
timestamp 1607639953
transform 1 0 56286 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1607639953
transform 1 0 57206 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_617
timestamp 1607639953
transform 1 0 57850 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_623
timestamp 1607639953
transform 1 0 58402 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1607639953
transform -1 0 58862 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1607639953
transform -1 0 58862 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1607639953
transform 1 0 2466 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1607639953
transform 1 0 1362 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1607639953
transform 1 0 1086 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1607639953
transform 1 0 4674 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1607639953
transform 1 0 3570 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_65
timestamp 1607639953
transform 1 0 7066 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1607639953
transform 1 0 6514 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1607639953
transform 1 0 5778 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1607639953
transform 1 0 6698 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _087_
timestamp 1607639953
transform 1 0 6790 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_80
timestamp 1607639953
transform 1 0 8446 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_73
timestamp 1607639953
transform 1 0 7802 0 1 13600
box -38 -48 314 592
use INVX2  INVX2
timestamp 1608122862
transform 1 0 8078 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_21_104
timestamp 1607639953
transform 1 0 10654 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_92
timestamp 1607639953
transform 1 0 9550 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1607639953
transform 1 0 12402 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_116
timestamp 1607639953
transform 1 0 11758 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1607639953
transform 1 0 12310 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1607639953
transform 1 0 14610 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1607639953
transform 1 0 13506 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1607639953
transform 1 0 16818 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1607639953
transform 1 0 15714 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1607639953
transform 1 0 19118 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1607639953
transform 1 0 18014 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1607639953
transform 1 0 17922 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1607639953
transform 1 0 21326 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1607639953
transform 1 0 20222 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_232
timestamp 1607639953
transform 1 0 22430 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1607639953
transform 1 0 24730 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1607639953
transform 1 0 23626 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1607639953
transform 1 0 23534 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_284
timestamp 1607639953
transform 1 0 27214 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_272
timestamp 1607639953
transform 1 0 26110 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _151_
timestamp 1607639953
transform 1 0 25834 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_306
timestamp 1607639953
transform 1 0 29238 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_304
timestamp 1607639953
transform 1 0 29054 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_296
timestamp 1607639953
transform 1 0 28318 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1607639953
transform 1 0 29146 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_330
timestamp 1607639953
transform 1 0 31446 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_318
timestamp 1607639953
transform 1 0 30342 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_342
timestamp 1607639953
transform 1 0 32550 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_367
timestamp 1607639953
transform 1 0 34850 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_354
timestamp 1607639953
transform 1 0 33654 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1607639953
transform 1 0 34758 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_391
timestamp 1607639953
transform 1 0 37058 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_379
timestamp 1607639953
transform 1 0 35954 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_415
timestamp 1607639953
transform 1 0 39266 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_403
timestamp 1607639953
transform 1 0 38162 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_440
timestamp 1607639953
transform 1 0 41566 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_428
timestamp 1607639953
transform 1 0 40462 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1607639953
transform 1 0 40370 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_452
timestamp 1607639953
transform 1 0 42670 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_476
timestamp 1607639953
transform 1 0 44878 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_464
timestamp 1607639953
transform 1 0 43774 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_501
timestamp 1607639953
transform 1 0 47178 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_489
timestamp 1607639953
transform 1 0 46074 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1607639953
transform 1 0 45982 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_525
timestamp 1607639953
transform 1 0 49386 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_513
timestamp 1607639953
transform 1 0 48282 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_550
timestamp 1607639953
transform 1 0 51686 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_545
timestamp 1607639953
transform 1 0 51226 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_533
timestamp 1607639953
transform 1 0 50122 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_529
timestamp 1607639953
transform 1 0 49754 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1607639953
transform 1 0 51594 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _010_
timestamp 1607639953
transform 1 0 49846 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_562
timestamp 1607639953
transform 1 0 52790 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_586
timestamp 1607639953
transform 1 0 54998 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_574
timestamp 1607639953
transform 1 0 53894 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_611
timestamp 1607639953
transform 1 0 57298 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_598
timestamp 1607639953
transform 1 0 56102 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1607639953
transform 1 0 57206 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_623
timestamp 1607639953
transform 1 0 58402 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1607639953
transform -1 0 58862 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1607639953
transform 1 0 2466 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1607639953
transform 1 0 1362 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1607639953
transform 1 0 1086 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1607639953
transform 1 0 5134 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1607639953
transform 1 0 4030 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1607639953
transform 1 0 3570 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1607639953
transform 1 0 3938 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1607639953
transform 1 0 6238 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1607639953
transform 1 0 8446 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1607639953
transform 1 0 7342 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1607639953
transform 1 0 10746 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1607639953
transform 1 0 9642 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1607639953
transform 1 0 9550 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1607639953
transform 1 0 12954 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1607639953
transform 1 0 11850 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1607639953
transform 1 0 15254 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1607639953
transform 1 0 14058 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1607639953
transform 1 0 15162 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1607639953
transform 1 0 16358 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1607639953
transform 1 0 18566 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1607639953
transform 1 0 17462 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1607639953
transform 1 0 20866 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1607639953
transform 1 0 19670 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1607639953
transform 1 0 20774 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1607639953
transform 1 0 23074 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1607639953
transform 1 0 21970 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_263
timestamp 1607639953
transform 1 0 25282 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_251
timestamp 1607639953
transform 1 0 24178 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_276
timestamp 1607639953
transform 1 0 26478 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_269
timestamp 1607639953
transform 1 0 25834 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1607639953
transform 1 0 26386 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _198_
timestamp 1607639953
transform 1 0 25558 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_300
timestamp 1607639953
transform 1 0 28686 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_288
timestamp 1607639953
transform 1 0 27582 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_324
timestamp 1607639953
transform 1 0 30894 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_320
timestamp 1607639953
transform 1 0 30526 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_312
timestamp 1607639953
transform 1 0 29790 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _192_
timestamp 1607639953
transform 1 0 30618 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_349
timestamp 1607639953
transform 1 0 33194 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_337
timestamp 1607639953
transform 1 0 32090 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1607639953
transform 1 0 31998 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_373
timestamp 1607639953
transform 1 0 35402 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_361
timestamp 1607639953
transform 1 0 34298 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_391
timestamp 1607639953
transform 1 0 37058 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_385
timestamp 1607639953
transform 1 0 36506 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _133_
timestamp 1607639953
transform 1 0 36782 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_410
timestamp 1607639953
transform 1 0 38806 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_398
timestamp 1607639953
transform 1 0 37702 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1607639953
transform 1 0 37610 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_434
timestamp 1607639953
transform 1 0 41014 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_422
timestamp 1607639953
transform 1 0 39910 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_459
timestamp 1607639953
transform 1 0 43314 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_446
timestamp 1607639953
transform 1 0 42118 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1607639953
transform 1 0 43222 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_474
timestamp 1607639953
transform 1 0 44694 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1607639953
transform 1 0 44418 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_498
timestamp 1607639953
transform 1 0 46902 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_486
timestamp 1607639953
transform 1 0 45798 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_520
timestamp 1607639953
transform 1 0 48926 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_518
timestamp 1607639953
transform 1 0 48742 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_510
timestamp 1607639953
transform 1 0 48006 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1607639953
transform 1 0 48834 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_544
timestamp 1607639953
transform 1 0 51134 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_532
timestamp 1607639953
transform 1 0 50030 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_565
timestamp 1607639953
transform 1 0 53066 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_556
timestamp 1607639953
transform 1 0 52238 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _152_
timestamp 1607639953
transform 1 0 52790 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_593
timestamp 1607639953
transform 1 0 55642 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_581
timestamp 1607639953
transform 1 0 54538 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_577
timestamp 1607639953
transform 1 0 54170 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1607639953
transform 1 0 54446 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_605
timestamp 1607639953
transform 1 0 56746 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_617
timestamp 1607639953
transform 1 0 57850 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1607639953
transform -1 0 58862 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1607639953
transform 1 0 2466 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1607639953
transform 1 0 1362 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1607639953
transform 1 0 1086 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_33
timestamp 1607639953
transform 1 0 4122 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_27
timestamp 1607639953
transform 1 0 3570 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _176_
timestamp 1607639953
transform 1 0 3846 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1607639953
transform 1 0 6790 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1607639953
transform 1 0 6330 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_45
timestamp 1607639953
transform 1 0 5226 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1607639953
transform 1 0 6698 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_82
timestamp 1607639953
transform 1 0 8630 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_74
timestamp 1607639953
transform 1 0 7894 0 1 14688
box -38 -48 222 592
use INVX4  INVX4
timestamp 1608122862
transform 1 0 8078 0 1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_23_106
timestamp 1607639953
transform 1 0 10838 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_94
timestamp 1607639953
transform 1 0 9734 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_131
timestamp 1607639953
transform 1 0 13138 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_127
timestamp 1607639953
transform 1 0 12770 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_123
timestamp 1607639953
transform 1 0 12402 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_118
timestamp 1607639953
transform 1 0 11942 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1607639953
transform 1 0 12310 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _208_
timestamp 1607639953
transform 1 0 12862 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_154
timestamp 1607639953
transform 1 0 15254 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_143
timestamp 1607639953
transform 1 0 14242 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _023_
timestamp 1607639953
transform 1 0 14978 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_166
timestamp 1607639953
transform 1 0 16358 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1607639953
transform 1 0 19118 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1607639953
transform 1 0 18014 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1607639953
transform 1 0 17830 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_178
timestamp 1607639953
transform 1 0 17462 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1607639953
transform 1 0 17922 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1607639953
transform 1 0 21326 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1607639953
transform 1 0 20222 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1607639953
transform 1 0 22430 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1607639953
transform 1 0 24730 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1607639953
transform 1 0 23626 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1607639953
transform 1 0 23534 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1607639953
transform 1 0 26938 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_269
timestamp 1607639953
transform 1 0 25834 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_306
timestamp 1607639953
transform 1 0 29238 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1607639953
transform 1 0 28042 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1607639953
transform 1 0 29146 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_328
timestamp 1607639953
transform 1 0 31262 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_324
timestamp 1607639953
transform 1 0 30894 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_318
timestamp 1607639953
transform 1 0 30342 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _088_
timestamp 1607639953
transform 1 0 30986 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_352
timestamp 1607639953
transform 1 0 33470 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_340
timestamp 1607639953
transform 1 0 32366 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_367
timestamp 1607639953
transform 1 0 34850 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_364
timestamp 1607639953
transform 1 0 34574 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1607639953
transform 1 0 34758 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_391
timestamp 1607639953
transform 1 0 37058 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_379
timestamp 1607639953
transform 1 0 35954 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_415
timestamp 1607639953
transform 1 0 39266 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_403
timestamp 1607639953
transform 1 0 38162 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_440
timestamp 1607639953
transform 1 0 41566 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_428
timestamp 1607639953
transform 1 0 40462 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1607639953
transform 1 0 40370 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_452
timestamp 1607639953
transform 1 0 42670 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_476
timestamp 1607639953
transform 1 0 44878 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_464
timestamp 1607639953
transform 1 0 43774 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_501
timestamp 1607639953
transform 1 0 47178 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_489
timestamp 1607639953
transform 1 0 46074 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1607639953
transform 1 0 45982 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_525
timestamp 1607639953
transform 1 0 49386 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_513
timestamp 1607639953
transform 1 0 48282 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_550
timestamp 1607639953
transform 1 0 51686 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_537
timestamp 1607639953
transform 1 0 50490 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1607639953
transform 1 0 51594 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_562
timestamp 1607639953
transform 1 0 52790 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_586
timestamp 1607639953
transform 1 0 54998 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_574
timestamp 1607639953
transform 1 0 53894 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_616
timestamp 1607639953
transform 1 0 57758 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_611
timestamp 1607639953
transform 1 0 57298 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_598
timestamp 1607639953
transform 1 0 56102 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1607639953
transform 1 0 57206 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _134_
timestamp 1607639953
transform 1 0 57482 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_624
timestamp 1607639953
transform 1 0 58494 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1607639953
transform -1 0 58862 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1607639953
transform 1 0 2466 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1607639953
transform 1 0 1362 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1607639953
transform 1 0 1086 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1607639953
transform 1 0 5134 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1607639953
transform 1 0 4030 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1607639953
transform 1 0 3570 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1607639953
transform 1 0 3938 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1607639953
transform 1 0 6238 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1607639953
transform 1 0 8446 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1607639953
transform 1 0 7342 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1607639953
transform 1 0 10746 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1607639953
transform 1 0 9642 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1607639953
transform 1 0 9550 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1607639953
transform 1 0 12954 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1607639953
transform 1 0 11850 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1607639953
transform 1 0 15254 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1607639953
transform 1 0 14058 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1607639953
transform 1 0 15162 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1607639953
transform 1 0 16358 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1607639953
transform 1 0 18566 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1607639953
transform 1 0 17462 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1607639953
transform 1 0 20866 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1607639953
transform 1 0 19670 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1607639953
transform 1 0 20774 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1607639953
transform 1 0 23074 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1607639953
transform 1 0 21970 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1607639953
transform 1 0 25282 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1607639953
transform 1 0 24178 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_279
timestamp 1607639953
transform 1 0 26754 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1607639953
transform 1 0 26386 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _168_
timestamp 1607639953
transform 1 0 26478 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_303
timestamp 1607639953
transform 1 0 28962 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_291
timestamp 1607639953
transform 1 0 27858 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_327
timestamp 1607639953
transform 1 0 31170 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_315
timestamp 1607639953
transform 1 0 30066 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_349
timestamp 1607639953
transform 1 0 33194 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_337
timestamp 1607639953
transform 1 0 32090 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_335
timestamp 1607639953
transform 1 0 31906 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1607639953
transform 1 0 31998 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_373
timestamp 1607639953
transform 1 0 35402 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_361
timestamp 1607639953
transform 1 0 34298 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_385
timestamp 1607639953
transform 1 0 36506 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_410
timestamp 1607639953
transform 1 0 38806 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_398
timestamp 1607639953
transform 1 0 37702 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1607639953
transform 1 0 37610 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_434
timestamp 1607639953
transform 1 0 41014 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_422
timestamp 1607639953
transform 1 0 39910 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_459
timestamp 1607639953
transform 1 0 43314 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_446
timestamp 1607639953
transform 1 0 42118 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1607639953
transform 1 0 43222 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_483
timestamp 1607639953
transform 1 0 45522 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_471
timestamp 1607639953
transform 1 0 44418 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_495
timestamp 1607639953
transform 1 0 46626 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_520
timestamp 1607639953
transform 1 0 48926 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_507
timestamp 1607639953
transform 1 0 47730 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1607639953
transform 1 0 48834 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_544
timestamp 1607639953
transform 1 0 51134 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_532
timestamp 1607639953
transform 1 0 50030 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_568
timestamp 1607639953
transform 1 0 53342 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_556
timestamp 1607639953
transform 1 0 52238 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_593
timestamp 1607639953
transform 1 0 55642 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_581
timestamp 1607639953
transform 1 0 54538 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1607639953
transform 1 0 54446 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1607639953
transform 1 0 55734 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_609
timestamp 1607639953
transform 1 0 57114 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_597
timestamp 1607639953
transform 1 0 56010 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_621
timestamp 1607639953
transform 1 0 58218 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1607639953
transform -1 0 58862 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_21
timestamp 1607639953
transform 1 0 3018 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_15
timestamp 1607639953
transform 1 0 2466 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1607639953
transform 1 0 1362 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1607639953
transform 1 0 1086 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _130_
timestamp 1607639953
transform 1 0 2742 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_33
timestamp 1607639953
transform 1 0 4122 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1607639953
transform 1 0 6790 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1607639953
transform 1 0 6330 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_45
timestamp 1607639953
transform 1 0 5226 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1607639953
transform 1 0 6698 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1607639953
transform 1 0 8998 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_74
timestamp 1607639953
transform 1 0 7894 0 1 15776
box -38 -48 222 592
use INVX8  INVX8
timestamp 1608122862
transform 1 0 8078 0 1 15776
box 0 -48 920 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1607639953
transform 1 0 11206 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1607639953
transform 1 0 10102 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1607639953
transform 1 0 12402 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1607639953
transform 1 0 12310 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1607639953
transform 1 0 14610 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1607639953
transform 1 0 13506 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1607639953
transform 1 0 16818 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1607639953
transform 1 0 15714 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1607639953
transform 1 0 19118 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1607639953
transform 1 0 18014 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1607639953
transform 1 0 17922 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1607639953
transform 1 0 21326 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1607639953
transform 1 0 20222 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1607639953
transform 1 0 22430 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1607639953
transform 1 0 24730 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1607639953
transform 1 0 23626 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1607639953
transform 1 0 23534 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_281
timestamp 1607639953
transform 1 0 26938 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_269
timestamp 1607639953
transform 1 0 25834 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_306
timestamp 1607639953
transform 1 0 29238 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_302
timestamp 1607639953
transform 1 0 28870 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_294
timestamp 1607639953
transform 1 0 28134 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_289
timestamp 1607639953
transform 1 0 27674 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1607639953
transform 1 0 29146 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _002_
timestamp 1607639953
transform 1 0 27858 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_330
timestamp 1607639953
transform 1 0 31446 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_318
timestamp 1607639953
transform 1 0 30342 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_344
timestamp 1607639953
transform 1 0 32734 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_338
timestamp 1607639953
transform 1 0 32182 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1607639953
transform 1 0 32458 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_370
timestamp 1607639953
transform 1 0 35126 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_365
timestamp 1607639953
transform 1 0 34666 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_356
timestamp 1607639953
transform 1 0 33838 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1607639953
transform 1 0 34758 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _143_
timestamp 1607639953
transform 1 0 34390 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _105_
timestamp 1607639953
transform 1 0 34850 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_394
timestamp 1607639953
transform 1 0 37334 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_382
timestamp 1607639953
transform 1 0 36230 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_418
timestamp 1607639953
transform 1 0 39542 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_406
timestamp 1607639953
transform 1 0 38438 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_440
timestamp 1607639953
transform 1 0 41566 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_428
timestamp 1607639953
transform 1 0 40462 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_426
timestamp 1607639953
transform 1 0 40278 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1607639953
transform 1 0 40370 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_452
timestamp 1607639953
transform 1 0 42670 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_476
timestamp 1607639953
transform 1 0 44878 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_464
timestamp 1607639953
transform 1 0 43774 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_501
timestamp 1607639953
transform 1 0 47178 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_489
timestamp 1607639953
transform 1 0 46074 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1607639953
transform 1 0 45982 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_525
timestamp 1607639953
transform 1 0 49386 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_513
timestamp 1607639953
transform 1 0 48282 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_550
timestamp 1607639953
transform 1 0 51686 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_537
timestamp 1607639953
transform 1 0 50490 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1607639953
transform 1 0 51594 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_562
timestamp 1607639953
transform 1 0 52790 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_586
timestamp 1607639953
transform 1 0 54998 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_574
timestamp 1607639953
transform 1 0 53894 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_611
timestamp 1607639953
transform 1 0 57298 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_598
timestamp 1607639953
transform 1 0 56102 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1607639953
transform 1 0 57206 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_623
timestamp 1607639953
transform 1 0 58402 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1607639953
transform -1 0 58862 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1607639953
transform 1 0 2466 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1607639953
transform 1 0 1362 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1607639953
transform 1 0 2466 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1607639953
transform 1 0 1362 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1607639953
transform 1 0 1086 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1607639953
transform 1 0 1086 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1607639953
transform 1 0 4674 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1607639953
transform 1 0 3570 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1607639953
transform 1 0 5134 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1607639953
transform 1 0 4030 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1607639953
transform 1 0 3570 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1607639953
transform 1 0 3938 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1607639953
transform 1 0 6790 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1607639953
transform 1 0 6514 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1607639953
transform 1 0 5778 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1607639953
transform 1 0 6238 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1607639953
transform 1 0 6698 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_74
timestamp 1607639953
transform 1 0 7894 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1607639953
transform 1 0 8446 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1607639953
transform 1 0 7342 0 -1 16864
box -38 -48 1142 592
use LATCH  LATCH
timestamp 1608122862
transform 1 0 8078 0 1 16864
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILLER_27_102
timestamp 1607639953
transform 1 0 10470 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_90
timestamp 1607639953
transform 1 0 9366 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1607639953
transform 1 0 10746 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1607639953
transform 1 0 9642 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1607639953
transform 1 0 9550 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1607639953
transform 1 0 12402 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_114
timestamp 1607639953
transform 1 0 11574 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1607639953
transform 1 0 12954 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1607639953
transform 1 0 11850 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1607639953
transform 1 0 12310 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1607639953
transform 1 0 14610 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1607639953
transform 1 0 13506 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1607639953
transform 1 0 15254 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1607639953
transform 1 0 14058 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1607639953
transform 1 0 15162 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1607639953
transform 1 0 16818 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1607639953
transform 1 0 15714 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1607639953
transform 1 0 16358 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1607639953
transform 1 0 19118 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1607639953
transform 1 0 18014 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1607639953
transform 1 0 18566 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1607639953
transform 1 0 17462 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1607639953
transform 1 0 17922 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1607639953
transform 1 0 21326 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1607639953
transform 1 0 20222 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1607639953
transform 1 0 20866 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1607639953
transform 1 0 19670 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1607639953
transform 1 0 20774 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1607639953
transform 1 0 22430 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1607639953
transform 1 0 23074 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1607639953
transform 1 0 21970 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1607639953
transform 1 0 24730 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1607639953
transform 1 0 23626 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1607639953
transform 1 0 25282 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1607639953
transform 1 0 24178 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1607639953
transform 1 0 23534 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1607639953
transform 1 0 26938 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_269
timestamp 1607639953
transform 1 0 25834 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_276
timestamp 1607639953
transform 1 0 26478 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1607639953
transform 1 0 26386 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_306
timestamp 1607639953
transform 1 0 29238 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1607639953
transform 1 0 28042 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_300
timestamp 1607639953
transform 1 0 28686 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_288
timestamp 1607639953
transform 1 0 27582 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1607639953
transform 1 0 29146 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_330
timestamp 1607639953
transform 1 0 31446 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_318
timestamp 1607639953
transform 1 0 30342 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_324
timestamp 1607639953
transform 1 0 30894 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_312
timestamp 1607639953
transform 1 0 29790 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_342
timestamp 1607639953
transform 1 0 32550 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_349
timestamp 1607639953
transform 1 0 33194 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_337
timestamp 1607639953
transform 1 0 32090 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1607639953
transform 1 0 31998 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_367
timestamp 1607639953
transform 1 0 34850 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_354
timestamp 1607639953
transform 1 0 33654 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_373
timestamp 1607639953
transform 1 0 35402 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_361
timestamp 1607639953
transform 1 0 34298 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1607639953
transform 1 0 34758 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_391
timestamp 1607639953
transform 1 0 37058 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_379
timestamp 1607639953
transform 1 0 35954 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_385
timestamp 1607639953
transform 1 0 36506 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_415
timestamp 1607639953
transform 1 0 39266 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_403
timestamp 1607639953
transform 1 0 38162 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_410
timestamp 1607639953
transform 1 0 38806 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_398
timestamp 1607639953
transform 1 0 37702 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1607639953
transform 1 0 37610 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_440
timestamp 1607639953
transform 1 0 41566 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_428
timestamp 1607639953
transform 1 0 40462 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_434
timestamp 1607639953
transform 1 0 41014 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_422
timestamp 1607639953
transform 1 0 39910 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1607639953
transform 1 0 40370 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_452
timestamp 1607639953
transform 1 0 42670 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_459
timestamp 1607639953
transform 1 0 43314 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_446
timestamp 1607639953
transform 1 0 42118 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1607639953
transform 1 0 43222 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_476
timestamp 1607639953
transform 1 0 44878 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_464
timestamp 1607639953
transform 1 0 43774 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_483
timestamp 1607639953
transform 1 0 45522 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_471
timestamp 1607639953
transform 1 0 44418 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_501
timestamp 1607639953
transform 1 0 47178 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_489
timestamp 1607639953
transform 1 0 46074 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_495
timestamp 1607639953
transform 1 0 46626 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1607639953
transform 1 0 45982 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_525
timestamp 1607639953
transform 1 0 49386 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_513
timestamp 1607639953
transform 1 0 48282 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_520
timestamp 1607639953
transform 1 0 48926 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_507
timestamp 1607639953
transform 1 0 47730 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1607639953
transform 1 0 48834 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_550
timestamp 1607639953
transform 1 0 51686 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_537
timestamp 1607639953
transform 1 0 50490 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_544
timestamp 1607639953
transform 1 0 51134 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_532
timestamp 1607639953
transform 1 0 50030 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1607639953
transform 1 0 51594 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_562
timestamp 1607639953
transform 1 0 52790 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_568
timestamp 1607639953
transform 1 0 53342 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_556
timestamp 1607639953
transform 1 0 52238 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_586
timestamp 1607639953
transform 1 0 54998 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_574
timestamp 1607639953
transform 1 0 53894 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_593
timestamp 1607639953
transform 1 0 55642 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_581
timestamp 1607639953
transform 1 0 54538 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1607639953
transform 1 0 54446 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_611
timestamp 1607639953
transform 1 0 57298 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_598
timestamp 1607639953
transform 1 0 56102 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_605
timestamp 1607639953
transform 1 0 56746 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1607639953
transform 1 0 57206 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_623
timestamp 1607639953
transform 1 0 58402 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_617
timestamp 1607639953
transform 1 0 57850 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1607639953
transform -1 0 58862 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1607639953
transform -1 0 58862 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1607639953
transform 1 0 2466 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1607639953
transform 1 0 1362 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1607639953
transform 1 0 1086 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1607639953
transform 1 0 5134 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1607639953
transform 1 0 4030 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1607639953
transform 1 0 3570 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1607639953
transform 1 0 3938 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1607639953
transform 1 0 6238 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_80
timestamp 1607639953
transform 1 0 8446 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1607639953
transform 1 0 7342 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _165_
timestamp 1607639953
transform 1 0 9182 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1607639953
transform 1 0 10746 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1607639953
transform 1 0 9642 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1607639953
transform 1 0 9458 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1607639953
transform 1 0 9550 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1607639953
transform 1 0 12954 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1607639953
transform 1 0 11850 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1607639953
transform 1 0 15254 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1607639953
transform 1 0 14058 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1607639953
transform 1 0 15162 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1607639953
transform 1 0 16358 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1607639953
transform 1 0 18566 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1607639953
transform 1 0 17462 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1607639953
transform 1 0 20866 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1607639953
transform 1 0 19670 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1607639953
transform 1 0 20774 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_239
timestamp 1607639953
transform 1 0 23074 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1607639953
transform 1 0 21970 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_264
timestamp 1607639953
transform 1 0 25374 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_252
timestamp 1607639953
transform 1 0 24270 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_247
timestamp 1607639953
transform 1 0 23810 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1607639953
transform 1 0 23994 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1607639953
transform 1 0 26478 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_272
timestamp 1607639953
transform 1 0 26110 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1607639953
transform 1 0 26386 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_300
timestamp 1607639953
transform 1 0 28686 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_288
timestamp 1607639953
transform 1 0 27582 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_324
timestamp 1607639953
transform 1 0 30894 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_312
timestamp 1607639953
transform 1 0 29790 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_349
timestamp 1607639953
transform 1 0 33194 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_337
timestamp 1607639953
transform 1 0 32090 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1607639953
transform 1 0 31998 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_361
timestamp 1607639953
transform 1 0 34298 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _014_
timestamp 1607639953
transform 1 0 35402 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_396
timestamp 1607639953
transform 1 0 37518 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_388
timestamp 1607639953
transform 1 0 36782 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_376
timestamp 1607639953
transform 1 0 35678 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_416
timestamp 1607639953
transform 1 0 39358 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_404
timestamp 1607639953
transform 1 0 38254 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_398
timestamp 1607639953
transform 1 0 37702 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1607639953
transform 1 0 37610 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _156_
timestamp 1607639953
transform 1 0 37978 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_440
timestamp 1607639953
transform 1 0 41566 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_428
timestamp 1607639953
transform 1 0 40462 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_459
timestamp 1607639953
transform 1 0 43314 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_452
timestamp 1607639953
transform 1 0 42670 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1607639953
transform 1 0 43222 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_483
timestamp 1607639953
transform 1 0 45522 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_471
timestamp 1607639953
transform 1 0 44418 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_495
timestamp 1607639953
transform 1 0 46626 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_520
timestamp 1607639953
transform 1 0 48926 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_507
timestamp 1607639953
transform 1 0 47730 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1607639953
transform 1 0 48834 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_544
timestamp 1607639953
transform 1 0 51134 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_532
timestamp 1607639953
transform 1 0 50030 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_568
timestamp 1607639953
transform 1 0 53342 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_556
timestamp 1607639953
transform 1 0 52238 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_593
timestamp 1607639953
transform 1 0 55642 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_581
timestamp 1607639953
transform 1 0 54538 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1607639953
transform 1 0 54446 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_605
timestamp 1607639953
transform 1 0 56746 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_617
timestamp 1607639953
transform 1 0 57850 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1607639953
transform -1 0 58862 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_17
timestamp 1607639953
transform 1 0 2650 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_11
timestamp 1607639953
transform 1 0 2098 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1607639953
transform 1 0 1362 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1607639953
transform 1 0 1086 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _068_
timestamp 1607639953
transform 1 0 2374 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_41
timestamp 1607639953
transform 1 0 4858 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_29
timestamp 1607639953
transform 1 0 3754 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1607639953
transform 1 0 6790 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_53
timestamp 1607639953
transform 1 0 5962 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1607639953
transform 1 0 6698 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_88
timestamp 1607639953
transform 1 0 9182 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_74
timestamp 1607639953
transform 1 0 7894 0 1 17952
box -38 -48 222 592
use MUX2X1  MUX2X1
timestamp 1608122862
transform 1 0 8078 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_29_100
timestamp 1607639953
transform 1 0 10286 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1607639953
transform 1 0 12402 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1607639953
transform 1 0 12126 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_112
timestamp 1607639953
transform 1 0 11390 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1607639953
transform 1 0 12310 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1607639953
transform 1 0 14610 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1607639953
transform 1 0 13506 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1607639953
transform 1 0 16818 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1607639953
transform 1 0 15714 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1607639953
transform 1 0 19118 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1607639953
transform 1 0 18014 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1607639953
transform 1 0 17922 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1607639953
transform 1 0 21326 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1607639953
transform 1 0 20222 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1607639953
transform 1 0 22430 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1607639953
transform 1 0 24730 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1607639953
transform 1 0 23626 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1607639953
transform 1 0 23534 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1607639953
transform 1 0 26938 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_269
timestamp 1607639953
transform 1 0 25834 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_306
timestamp 1607639953
transform 1 0 29238 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1607639953
transform 1 0 28042 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1607639953
transform 1 0 29146 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_330
timestamp 1607639953
transform 1 0 31446 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_318
timestamp 1607639953
transform 1 0 30342 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_342
timestamp 1607639953
transform 1 0 32550 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_367
timestamp 1607639953
transform 1 0 34850 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_354
timestamp 1607639953
transform 1 0 33654 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1607639953
transform 1 0 34758 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_391
timestamp 1607639953
transform 1 0 37058 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_379
timestamp 1607639953
transform 1 0 35954 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_415
timestamp 1607639953
transform 1 0 39266 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_403
timestamp 1607639953
transform 1 0 38162 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_440
timestamp 1607639953
transform 1 0 41566 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_428
timestamp 1607639953
transform 1 0 40462 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1607639953
transform 1 0 40370 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_452
timestamp 1607639953
transform 1 0 42670 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_476
timestamp 1607639953
transform 1 0 44878 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_464
timestamp 1607639953
transform 1 0 43774 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_501
timestamp 1607639953
transform 1 0 47178 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_497
timestamp 1607639953
transform 1 0 46810 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_489
timestamp 1607639953
transform 1 0 46074 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1607639953
transform 1 0 45982 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _171_
timestamp 1607639953
transform 1 0 46902 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_525
timestamp 1607639953
transform 1 0 49386 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_513
timestamp 1607639953
transform 1 0 48282 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_550
timestamp 1607639953
transform 1 0 51686 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_537
timestamp 1607639953
transform 1 0 50490 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1607639953
transform 1 0 51594 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_570
timestamp 1607639953
transform 1 0 53526 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_562
timestamp 1607639953
transform 1 0 52790 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_588
timestamp 1607639953
transform 1 0 55182 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_576
timestamp 1607639953
transform 1 0 54078 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _119_
timestamp 1607639953
transform 1 0 53802 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_611
timestamp 1607639953
transform 1 0 57298 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_608
timestamp 1607639953
transform 1 0 57022 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_600
timestamp 1607639953
transform 1 0 56286 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1607639953
transform 1 0 57206 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_623
timestamp 1607639953
transform 1 0 58402 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1607639953
transform -1 0 58862 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1607639953
transform 1 0 2466 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1607639953
transform 1 0 1362 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1607639953
transform 1 0 1086 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1607639953
transform 1 0 5134 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1607639953
transform 1 0 4030 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1607639953
transform 1 0 3570 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1607639953
transform 1 0 3938 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1607639953
transform 1 0 6238 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1607639953
transform 1 0 8446 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1607639953
transform 1 0 7342 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1607639953
transform 1 0 10746 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1607639953
transform 1 0 9642 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1607639953
transform 1 0 9550 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1607639953
transform 1 0 12954 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1607639953
transform 1 0 11850 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1607639953
transform 1 0 15254 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1607639953
transform 1 0 14058 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1607639953
transform 1 0 15162 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1607639953
transform 1 0 16358 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1607639953
transform 1 0 18566 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1607639953
transform 1 0 17462 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1607639953
transform 1 0 20866 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1607639953
transform 1 0 19670 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1607639953
transform 1 0 20774 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1607639953
transform 1 0 23074 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1607639953
transform 1 0 21970 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1607639953
transform 1 0 25282 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1607639953
transform 1 0 24178 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_276
timestamp 1607639953
transform 1 0 26478 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1607639953
transform 1 0 26386 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_300
timestamp 1607639953
transform 1 0 28686 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_288
timestamp 1607639953
transform 1 0 27582 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_324
timestamp 1607639953
transform 1 0 30894 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_312
timestamp 1607639953
transform 1 0 29790 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_349
timestamp 1607639953
transform 1 0 33194 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_337
timestamp 1607639953
transform 1 0 32090 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1607639953
transform 1 0 31998 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_371
timestamp 1607639953
transform 1 0 35218 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_367
timestamp 1607639953
transform 1 0 34850 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_361
timestamp 1607639953
transform 1 0 34298 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _175_
timestamp 1607639953
transform 1 0 34942 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_395
timestamp 1607639953
transform 1 0 37426 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_383
timestamp 1607639953
transform 1 0 36322 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_410
timestamp 1607639953
transform 1 0 38806 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_398
timestamp 1607639953
transform 1 0 37702 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1607639953
transform 1 0 37610 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_434
timestamp 1607639953
transform 1 0 41014 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_422
timestamp 1607639953
transform 1 0 39910 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_459
timestamp 1607639953
transform 1 0 43314 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_446
timestamp 1607639953
transform 1 0 42118 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1607639953
transform 1 0 43222 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_478
timestamp 1607639953
transform 1 0 45062 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_471
timestamp 1607639953
transform 1 0 44418 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _148_
timestamp 1607639953
transform 1 0 44786 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_502
timestamp 1607639953
transform 1 0 47270 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_490
timestamp 1607639953
transform 1 0 46166 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_520
timestamp 1607639953
transform 1 0 48926 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_518
timestamp 1607639953
transform 1 0 48742 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_514
timestamp 1607639953
transform 1 0 48374 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1607639953
transform 1 0 48834 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_544
timestamp 1607639953
transform 1 0 51134 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_532
timestamp 1607639953
transform 1 0 50030 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_568
timestamp 1607639953
transform 1 0 53342 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_556
timestamp 1607639953
transform 1 0 52238 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_593
timestamp 1607639953
transform 1 0 55642 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_581
timestamp 1607639953
transform 1 0 54538 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1607639953
transform 1 0 54446 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_605
timestamp 1607639953
transform 1 0 56746 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_617
timestamp 1607639953
transform 1 0 57850 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1607639953
transform -1 0 58862 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1607639953
transform 1 0 2466 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1607639953
transform 1 0 1362 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1607639953
transform 1 0 1086 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_39
timestamp 1607639953
transform 1 0 4674 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1607639953
transform 1 0 3570 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_66
timestamp 1607639953
transform 1 0 7158 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_62
timestamp 1607639953
transform 1 0 6790 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_58
timestamp 1607639953
transform 1 0 6422 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_50
timestamp 1607639953
transform 1 0 5686 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1607639953
transform 1 0 6698 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _166_
timestamp 1607639953
transform 1 0 5410 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_82
timestamp 1607639953
transform 1 0 8630 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_70
timestamp 1607639953
transform 1 0 7526 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _022_
timestamp 1607639953
transform 1 0 7250 0 1 19040
box -38 -48 314 592
use NAND2X1  NAND2X1
timestamp 1608122862
transform 1 0 8078 0 1 19040
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_31_106
timestamp 1607639953
transform 1 0 10838 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_94
timestamp 1607639953
transform 1 0 9734 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1607639953
transform 1 0 12402 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_118
timestamp 1607639953
transform 1 0 11942 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1607639953
transform 1 0 12310 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1607639953
transform 1 0 14610 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1607639953
transform 1 0 13506 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1607639953
transform 1 0 16818 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1607639953
transform 1 0 15714 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1607639953
transform 1 0 19118 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1607639953
transform 1 0 18014 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1607639953
transform 1 0 17922 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1607639953
transform 1 0 21326 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1607639953
transform 1 0 20222 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1607639953
transform 1 0 22430 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1607639953
transform 1 0 24730 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1607639953
transform 1 0 23626 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1607639953
transform 1 0 23534 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1607639953
transform 1 0 26938 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_269
timestamp 1607639953
transform 1 0 25834 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_306
timestamp 1607639953
transform 1 0 29238 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1607639953
transform 1 0 28042 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1607639953
transform 1 0 29146 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_330
timestamp 1607639953
transform 1 0 31446 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_318
timestamp 1607639953
transform 1 0 30342 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_342
timestamp 1607639953
transform 1 0 32550 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_367
timestamp 1607639953
transform 1 0 34850 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_354
timestamp 1607639953
transform 1 0 33654 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1607639953
transform 1 0 34758 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_391
timestamp 1607639953
transform 1 0 37058 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_379
timestamp 1607639953
transform 1 0 35954 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_415
timestamp 1607639953
transform 1 0 39266 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_403
timestamp 1607639953
transform 1 0 38162 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_440
timestamp 1607639953
transform 1 0 41566 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_428
timestamp 1607639953
transform 1 0 40462 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1607639953
transform 1 0 40370 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_452
timestamp 1607639953
transform 1 0 42670 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_476
timestamp 1607639953
transform 1 0 44878 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_464
timestamp 1607639953
transform 1 0 43774 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_501
timestamp 1607639953
transform 1 0 47178 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_489
timestamp 1607639953
transform 1 0 46074 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1607639953
transform 1 0 45982 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_525
timestamp 1607639953
transform 1 0 49386 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_513
timestamp 1607639953
transform 1 0 48282 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_550
timestamp 1607639953
transform 1 0 51686 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_537
timestamp 1607639953
transform 1 0 50490 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1607639953
transform 1 0 51594 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_562
timestamp 1607639953
transform 1 0 52790 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_586
timestamp 1607639953
transform 1 0 54998 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_574
timestamp 1607639953
transform 1 0 53894 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_611
timestamp 1607639953
transform 1 0 57298 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_598
timestamp 1607639953
transform 1 0 56102 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1607639953
transform 1 0 57206 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_623
timestamp 1607639953
transform 1 0 58402 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1607639953
transform -1 0 58862 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1607639953
transform 1 0 2466 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1607639953
transform 1 0 1362 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1607639953
transform 1 0 1086 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1607639953
transform 1 0 5134 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1607639953
transform 1 0 4030 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1607639953
transform 1 0 3570 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1607639953
transform 1 0 3938 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1607639953
transform 1 0 6238 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1607639953
transform 1 0 8446 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1607639953
transform 1 0 7342 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1607639953
transform 1 0 10746 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1607639953
transform 1 0 9642 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1607639953
transform 1 0 9550 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1607639953
transform 1 0 12954 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1607639953
transform 1 0 11850 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1607639953
transform 1 0 15254 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1607639953
transform 1 0 14058 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1607639953
transform 1 0 15162 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1607639953
transform 1 0 16358 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1607639953
transform 1 0 18566 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1607639953
transform 1 0 17462 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1607639953
transform 1 0 20866 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1607639953
transform 1 0 19670 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1607639953
transform 1 0 20774 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1607639953
transform 1 0 23074 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1607639953
transform 1 0 21970 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1607639953
transform 1 0 25282 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1607639953
transform 1 0 24178 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_276
timestamp 1607639953
transform 1 0 26478 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1607639953
transform 1 0 26386 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_300
timestamp 1607639953
transform 1 0 28686 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_288
timestamp 1607639953
transform 1 0 27582 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_324
timestamp 1607639953
transform 1 0 30894 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_312
timestamp 1607639953
transform 1 0 29790 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_349
timestamp 1607639953
transform 1 0 33194 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_337
timestamp 1607639953
transform 1 0 32090 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1607639953
transform 1 0 31998 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_373
timestamp 1607639953
transform 1 0 35402 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_361
timestamp 1607639953
transform 1 0 34298 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_385
timestamp 1607639953
transform 1 0 36506 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_410
timestamp 1607639953
transform 1 0 38806 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_398
timestamp 1607639953
transform 1 0 37702 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1607639953
transform 1 0 37610 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_439
timestamp 1607639953
transform 1 0 41474 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_427
timestamp 1607639953
transform 1 0 40370 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_422
timestamp 1607639953
transform 1 0 39910 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1607639953
transform 1 0 40094 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_459
timestamp 1607639953
transform 1 0 43314 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_456
timestamp 1607639953
transform 1 0 43038 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_448
timestamp 1607639953
transform 1 0 42302 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1607639953
transform 1 0 43222 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1607639953
transform 1 0 42026 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_483
timestamp 1607639953
transform 1 0 45522 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_471
timestamp 1607639953
transform 1 0 44418 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_495
timestamp 1607639953
transform 1 0 46626 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_520
timestamp 1607639953
transform 1 0 48926 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_507
timestamp 1607639953
transform 1 0 47730 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1607639953
transform 1 0 48834 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_544
timestamp 1607639953
transform 1 0 51134 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_532
timestamp 1607639953
transform 1 0 50030 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_568
timestamp 1607639953
transform 1 0 53342 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_556
timestamp 1607639953
transform 1 0 52238 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_593
timestamp 1607639953
transform 1 0 55642 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_581
timestamp 1607639953
transform 1 0 54538 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1607639953
transform 1 0 54446 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_605
timestamp 1607639953
transform 1 0 56746 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_617
timestamp 1607639953
transform 1 0 57850 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1607639953
transform -1 0 58862 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1607639953
transform 1 0 2466 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1607639953
transform 1 0 1362 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1607639953
transform 1 0 2466 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1607639953
transform 1 0 1362 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1607639953
transform 1 0 1086 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1607639953
transform 1 0 1086 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1607639953
transform 1 0 5134 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1607639953
transform 1 0 4030 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1607639953
transform 1 0 3570 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1607639953
transform 1 0 4674 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1607639953
transform 1 0 3570 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1607639953
transform 1 0 3938 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1607639953
transform 1 0 6238 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1607639953
transform 1 0 6790 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1607639953
transform 1 0 6514 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1607639953
transform 1 0 5778 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1607639953
transform 1 0 6698 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1607639953
transform 1 0 8446 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1607639953
transform 1 0 7342 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_84
timestamp 1607639953
transform 1 0 8814 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_74
timestamp 1607639953
transform 1 0 7894 0 1 20128
box -38 -48 222 592
use NAND3X1  NAND3X1
timestamp 1608122862
transform 1 0 8078 0 1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1607639953
transform 1 0 10746 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1607639953
transform 1 0 9642 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_107
timestamp 1607639953
transform 1 0 10930 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_96
timestamp 1607639953
transform 1 0 9918 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1607639953
transform 1 0 9550 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _121_
timestamp 1607639953
transform 1 0 10654 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1607639953
transform 1 0 12954 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1607639953
transform 1 0 11850 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1607639953
transform 1 0 12402 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_119
timestamp 1607639953
transform 1 0 12034 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1607639953
transform 1 0 12310 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1607639953
transform 1 0 15254 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1607639953
transform 1 0 14058 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1607639953
transform 1 0 14610 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1607639953
transform 1 0 13506 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1607639953
transform 1 0 15162 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1607639953
transform 1 0 16358 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_171
timestamp 1607639953
transform 1 0 16818 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_159
timestamp 1607639953
transform 1 0 15714 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1607639953
transform 1 0 18566 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1607639953
transform 1 0 17462 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1607639953
transform 1 0 19118 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1607639953
transform 1 0 18014 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1607639953
transform 1 0 17922 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1607639953
transform 1 0 20866 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1607639953
transform 1 0 19670 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1607639953
transform 1 0 21326 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1607639953
transform 1 0 20222 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1607639953
transform 1 0 20774 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1607639953
transform 1 0 23074 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1607639953
transform 1 0 21970 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1607639953
transform 1 0 22430 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1607639953
transform 1 0 25282 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1607639953
transform 1 0 24178 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1607639953
transform 1 0 24730 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1607639953
transform 1 0 23626 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1607639953
transform 1 0 23534 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1607639953
transform 1 0 26478 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1607639953
transform 1 0 26938 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_269
timestamp 1607639953
transform 1 0 25834 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1607639953
transform 1 0 26386 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_300
timestamp 1607639953
transform 1 0 28686 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_288
timestamp 1607639953
transform 1 0 27582 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_306
timestamp 1607639953
transform 1 0 29238 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1607639953
transform 1 0 28042 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1607639953
transform 1 0 29146 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_324
timestamp 1607639953
transform 1 0 30894 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_312
timestamp 1607639953
transform 1 0 29790 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_330
timestamp 1607639953
transform 1 0 31446 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_318
timestamp 1607639953
transform 1 0 30342 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_349
timestamp 1607639953
transform 1 0 33194 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_337
timestamp 1607639953
transform 1 0 32090 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_342
timestamp 1607639953
transform 1 0 32550 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1607639953
transform 1 0 31998 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_373
timestamp 1607639953
transform 1 0 35402 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_361
timestamp 1607639953
transform 1 0 34298 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_367
timestamp 1607639953
transform 1 0 34850 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_354
timestamp 1607639953
transform 1 0 33654 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1607639953
transform 1 0 34758 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_385
timestamp 1607639953
transform 1 0 36506 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_391
timestamp 1607639953
transform 1 0 37058 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_379
timestamp 1607639953
transform 1 0 35954 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_410
timestamp 1607639953
transform 1 0 38806 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_398
timestamp 1607639953
transform 1 0 37702 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_415
timestamp 1607639953
transform 1 0 39266 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_403
timestamp 1607639953
transform 1 0 38162 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1607639953
transform 1 0 37610 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_434
timestamp 1607639953
transform 1 0 41014 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_422
timestamp 1607639953
transform 1 0 39910 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_440
timestamp 1607639953
transform 1 0 41566 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_428
timestamp 1607639953
transform 1 0 40462 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1607639953
transform 1 0 40370 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_459
timestamp 1607639953
transform 1 0 43314 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_446
timestamp 1607639953
transform 1 0 42118 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_452
timestamp 1607639953
transform 1 0 42670 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1607639953
transform 1 0 43222 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_483
timestamp 1607639953
transform 1 0 45522 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_471
timestamp 1607639953
transform 1 0 44418 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_476
timestamp 1607639953
transform 1 0 44878 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_464
timestamp 1607639953
transform 1 0 43774 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_495
timestamp 1607639953
transform 1 0 46626 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_501
timestamp 1607639953
transform 1 0 47178 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_489
timestamp 1607639953
transform 1 0 46074 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1607639953
transform 1 0 45982 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_520
timestamp 1607639953
transform 1 0 48926 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_507
timestamp 1607639953
transform 1 0 47730 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_525
timestamp 1607639953
transform 1 0 49386 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_513
timestamp 1607639953
transform 1 0 48282 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1607639953
transform 1 0 48834 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_544
timestamp 1607639953
transform 1 0 51134 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_532
timestamp 1607639953
transform 1 0 50030 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_550
timestamp 1607639953
transform 1 0 51686 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_537
timestamp 1607639953
transform 1 0 50490 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1607639953
transform 1 0 51594 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_568
timestamp 1607639953
transform 1 0 53342 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_556
timestamp 1607639953
transform 1 0 52238 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_562
timestamp 1607639953
transform 1 0 52790 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_593
timestamp 1607639953
transform 1 0 55642 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_581
timestamp 1607639953
transform 1 0 54538 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_586
timestamp 1607639953
transform 1 0 54998 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_574
timestamp 1607639953
transform 1 0 53894 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1607639953
transform 1 0 54446 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_605
timestamp 1607639953
transform 1 0 56746 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_611
timestamp 1607639953
transform 1 0 57298 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_609
timestamp 1607639953
transform 1 0 57114 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_603
timestamp 1607639953
transform 1 0 56562 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_598
timestamp 1607639953
transform 1 0 56102 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1607639953
transform 1 0 57206 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _195_
timestamp 1607639953
transform 1 0 56286 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_617
timestamp 1607639953
transform 1 0 57850 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_623
timestamp 1607639953
transform 1 0 58402 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1607639953
transform -1 0 58862 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1607639953
transform -1 0 58862 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1607639953
transform 1 0 2466 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1607639953
transform 1 0 1362 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1607639953
transform 1 0 1086 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1607639953
transform 1 0 4674 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1607639953
transform 1 0 3570 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1607639953
transform 1 0 6790 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1607639953
transform 1 0 6514 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1607639953
transform 1 0 5778 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1607639953
transform 1 0 6698 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_82
timestamp 1607639953
transform 1 0 8630 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_74
timestamp 1607639953
transform 1 0 7894 0 1 21216
box -38 -48 222 592
use NOR2X1  NOR2X1
timestamp 1608122862
transform 1 0 8078 0 1 21216
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_35_106
timestamp 1607639953
transform 1 0 10838 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1607639953
transform 1 0 9734 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1607639953
transform 1 0 12402 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_118
timestamp 1607639953
transform 1 0 11942 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1607639953
transform 1 0 12310 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_147
timestamp 1607639953
transform 1 0 14610 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_135
timestamp 1607639953
transform 1 0 13506 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_171
timestamp 1607639953
transform 1 0 16818 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_159
timestamp 1607639953
transform 1 0 15714 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1607639953
transform 1 0 19118 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1607639953
transform 1 0 18014 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1607639953
transform 1 0 17922 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1607639953
transform 1 0 21326 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1607639953
transform 1 0 20222 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1607639953
transform 1 0 22430 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1607639953
transform 1 0 24730 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1607639953
transform 1 0 23626 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1607639953
transform 1 0 23534 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1607639953
transform 1 0 26938 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_269
timestamp 1607639953
transform 1 0 25834 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_306
timestamp 1607639953
transform 1 0 29238 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1607639953
transform 1 0 28042 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1607639953
transform 1 0 29146 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_319
timestamp 1607639953
transform 1 0 30434 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_314
timestamp 1607639953
transform 1 0 29974 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _147_
timestamp 1607639953
transform 1 0 30158 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_343
timestamp 1607639953
transform 1 0 32642 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_331
timestamp 1607639953
transform 1 0 31538 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_367
timestamp 1607639953
transform 1 0 34850 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_363
timestamp 1607639953
transform 1 0 34482 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_355
timestamp 1607639953
transform 1 0 33746 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1607639953
transform 1 0 34758 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_391
timestamp 1607639953
transform 1 0 37058 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_379
timestamp 1607639953
transform 1 0 35954 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_415
timestamp 1607639953
transform 1 0 39266 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_403
timestamp 1607639953
transform 1 0 38162 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_440
timestamp 1607639953
transform 1 0 41566 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_428
timestamp 1607639953
transform 1 0 40462 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1607639953
transform 1 0 40370 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_452
timestamp 1607639953
transform 1 0 42670 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_476
timestamp 1607639953
transform 1 0 44878 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_464
timestamp 1607639953
transform 1 0 43774 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_501
timestamp 1607639953
transform 1 0 47178 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_489
timestamp 1607639953
transform 1 0 46074 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1607639953
transform 1 0 45982 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_525
timestamp 1607639953
transform 1 0 49386 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_513
timestamp 1607639953
transform 1 0 48282 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_550
timestamp 1607639953
transform 1 0 51686 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_537
timestamp 1607639953
transform 1 0 50490 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1607639953
transform 1 0 51594 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_562
timestamp 1607639953
transform 1 0 52790 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_586
timestamp 1607639953
transform 1 0 54998 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_574
timestamp 1607639953
transform 1 0 53894 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_611
timestamp 1607639953
transform 1 0 57298 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_598
timestamp 1607639953
transform 1 0 56102 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1607639953
transform 1 0 57206 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_623
timestamp 1607639953
transform 1 0 58402 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1607639953
transform -1 0 58862 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_22
timestamp 1607639953
transform 1 0 3110 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_15
timestamp 1607639953
transform 1 0 2466 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1607639953
transform 1 0 1362 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1607639953
transform 1 0 1086 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _011_
timestamp 1607639953
transform 1 0 2834 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1607639953
transform 1 0 5134 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1607639953
transform 1 0 4030 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_30
timestamp 1607639953
transform 1 0 3846 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1607639953
transform 1 0 3938 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1607639953
transform 1 0 6238 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1607639953
transform 1 0 8446 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1607639953
transform 1 0 7342 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1607639953
transform 1 0 10746 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1607639953
transform 1 0 9642 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1607639953
transform 1 0 9550 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1607639953
transform 1 0 12954 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_117
timestamp 1607639953
transform 1 0 11850 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1607639953
transform 1 0 15254 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1607639953
transform 1 0 14058 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1607639953
transform 1 0 15162 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_166
timestamp 1607639953
transform 1 0 16358 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_193
timestamp 1607639953
transform 1 0 18842 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_181
timestamp 1607639953
transform 1 0 17738 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1607639953
transform 1 0 17462 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_218
timestamp 1607639953
transform 1 0 21142 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1607639953
transform 1 0 20682 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_205
timestamp 1607639953
transform 1 0 19946 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1607639953
transform 1 0 20774 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1607639953
transform 1 0 20866 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_242
timestamp 1607639953
transform 1 0 23350 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_230
timestamp 1607639953
transform 1 0 22246 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_254
timestamp 1607639953
transform 1 0 24454 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_276
timestamp 1607639953
transform 1 0 26478 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_274
timestamp 1607639953
transform 1 0 26294 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_266
timestamp 1607639953
transform 1 0 25558 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1607639953
transform 1 0 26386 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_300
timestamp 1607639953
transform 1 0 28686 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_288
timestamp 1607639953
transform 1 0 27582 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_324
timestamp 1607639953
transform 1 0 30894 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_312
timestamp 1607639953
transform 1 0 29790 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_349
timestamp 1607639953
transform 1 0 33194 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_337
timestamp 1607639953
transform 1 0 32090 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1607639953
transform 1 0 31998 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_373
timestamp 1607639953
transform 1 0 35402 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_361
timestamp 1607639953
transform 1 0 34298 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_385
timestamp 1607639953
transform 1 0 36506 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_410
timestamp 1607639953
transform 1 0 38806 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_398
timestamp 1607639953
transform 1 0 37702 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1607639953
transform 1 0 37610 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_434
timestamp 1607639953
transform 1 0 41014 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_422
timestamp 1607639953
transform 1 0 39910 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_459
timestamp 1607639953
transform 1 0 43314 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_446
timestamp 1607639953
transform 1 0 42118 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1607639953
transform 1 0 43222 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_483
timestamp 1607639953
transform 1 0 45522 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_471
timestamp 1607639953
transform 1 0 44418 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_506
timestamp 1607639953
transform 1 0 47638 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_498
timestamp 1607639953
transform 1 0 46902 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _170_
timestamp 1607639953
transform 1 0 46626 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_520
timestamp 1607639953
transform 1 0 48926 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_518
timestamp 1607639953
transform 1 0 48742 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_510
timestamp 1607639953
transform 1 0 48006 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1607639953
transform 1 0 48834 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _149_
timestamp 1607639953
transform 1 0 47730 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_544
timestamp 1607639953
transform 1 0 51134 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_532
timestamp 1607639953
transform 1 0 50030 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_568
timestamp 1607639953
transform 1 0 53342 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_556
timestamp 1607639953
transform 1 0 52238 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_593
timestamp 1607639953
transform 1 0 55642 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_581
timestamp 1607639953
transform 1 0 54538 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1607639953
transform 1 0 54446 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_605
timestamp 1607639953
transform 1 0 56746 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_617
timestamp 1607639953
transform 1 0 57850 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1607639953
transform -1 0 58862 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1607639953
transform 1 0 2466 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1607639953
transform 1 0 1362 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1607639953
transform 1 0 1086 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1607639953
transform 1 0 4674 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1607639953
transform 1 0 3570 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1607639953
transform 1 0 6790 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1607639953
transform 1 0 6514 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1607639953
transform 1 0 5778 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1607639953
transform 1 0 6698 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_74
timestamp 1607639953
transform 1 0 7894 0 1 22304
box -38 -48 222 592
use NOR3X1  NOR3X1
timestamp 1608122862
transform 1 0 8078 0 1 22304
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILLER_37_102
timestamp 1607639953
transform 1 0 10470 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_90
timestamp 1607639953
transform 1 0 9366 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1607639953
transform 1 0 12402 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_114
timestamp 1607639953
transform 1 0 11574 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1607639953
transform 1 0 12310 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_147
timestamp 1607639953
transform 1 0 14610 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_135
timestamp 1607639953
transform 1 0 13506 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_171
timestamp 1607639953
transform 1 0 16818 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_159
timestamp 1607639953
transform 1 0 15714 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1607639953
transform 1 0 19118 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1607639953
transform 1 0 18014 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1607639953
transform 1 0 17922 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_220
timestamp 1607639953
transform 1 0 21326 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1607639953
transform 1 0 20222 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_232
timestamp 1607639953
transform 1 0 22430 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1607639953
transform 1 0 24730 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1607639953
transform 1 0 23626 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1607639953
transform 1 0 23534 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1607639953
transform 1 0 26938 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_269
timestamp 1607639953
transform 1 0 25834 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_306
timestamp 1607639953
transform 1 0 29238 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1607639953
transform 1 0 28042 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1607639953
transform 1 0 29146 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_330
timestamp 1607639953
transform 1 0 31446 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_318
timestamp 1607639953
transform 1 0 30342 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_342
timestamp 1607639953
transform 1 0 32550 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_367
timestamp 1607639953
transform 1 0 34850 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_354
timestamp 1607639953
transform 1 0 33654 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1607639953
transform 1 0 34758 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_394
timestamp 1607639953
transform 1 0 37334 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_382
timestamp 1607639953
transform 1 0 36230 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _083_
timestamp 1607639953
transform 1 0 35954 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_418
timestamp 1607639953
transform 1 0 39542 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_406
timestamp 1607639953
transform 1 0 38438 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_440
timestamp 1607639953
transform 1 0 41566 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_428
timestamp 1607639953
transform 1 0 40462 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_426
timestamp 1607639953
transform 1 0 40278 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1607639953
transform 1 0 40370 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_452
timestamp 1607639953
transform 1 0 42670 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_476
timestamp 1607639953
transform 1 0 44878 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_464
timestamp 1607639953
transform 1 0 43774 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_501
timestamp 1607639953
transform 1 0 47178 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_489
timestamp 1607639953
transform 1 0 46074 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1607639953
transform 1 0 45982 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_525
timestamp 1607639953
transform 1 0 49386 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_513
timestamp 1607639953
transform 1 0 48282 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_550
timestamp 1607639953
transform 1 0 51686 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_537
timestamp 1607639953
transform 1 0 50490 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1607639953
transform 1 0 51594 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_562
timestamp 1607639953
transform 1 0 52790 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_586
timestamp 1607639953
transform 1 0 54998 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_574
timestamp 1607639953
transform 1 0 53894 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _026_
timestamp 1607639953
transform 1 0 55734 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_611
timestamp 1607639953
transform 1 0 57298 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_609
timestamp 1607639953
transform 1 0 57114 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_597
timestamp 1607639953
transform 1 0 56010 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1607639953
transform 1 0 57206 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_623
timestamp 1607639953
transform 1 0 58402 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1607639953
transform -1 0 58862 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1607639953
transform 1 0 2466 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1607639953
transform 1 0 1362 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1607639953
transform 1 0 1086 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1607639953
transform 1 0 5134 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1607639953
transform 1 0 4030 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1607639953
transform 1 0 3570 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1607639953
transform 1 0 3938 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1607639953
transform 1 0 6238 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1607639953
transform 1 0 8446 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1607639953
transform 1 0 7342 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1607639953
transform 1 0 10746 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1607639953
transform 1 0 9642 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1607639953
transform 1 0 9550 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_129
timestamp 1607639953
transform 1 0 12954 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_117
timestamp 1607639953
transform 1 0 11850 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1607639953
transform 1 0 15254 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1607639953
transform 1 0 14058 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1607639953
transform 1 0 15162 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1607639953
transform 1 0 16358 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_190
timestamp 1607639953
transform 1 0 18566 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_178
timestamp 1607639953
transform 1 0 17462 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1607639953
transform 1 0 20866 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_202
timestamp 1607639953
transform 1 0 19670 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1607639953
transform 1 0 20774 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1607639953
transform 1 0 23074 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1607639953
transform 1 0 21970 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_263
timestamp 1607639953
transform 1 0 25282 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_251
timestamp 1607639953
transform 1 0 24178 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_276
timestamp 1607639953
transform 1 0 26478 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1607639953
transform 1 0 26386 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_300
timestamp 1607639953
transform 1 0 28686 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_288
timestamp 1607639953
transform 1 0 27582 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_324
timestamp 1607639953
transform 1 0 30894 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_312
timestamp 1607639953
transform 1 0 29790 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_349
timestamp 1607639953
transform 1 0 33194 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_337
timestamp 1607639953
transform 1 0 32090 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1607639953
transform 1 0 31998 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_373
timestamp 1607639953
transform 1 0 35402 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_361
timestamp 1607639953
transform 1 0 34298 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_385
timestamp 1607639953
transform 1 0 36506 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_410
timestamp 1607639953
transform 1 0 38806 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_398
timestamp 1607639953
transform 1 0 37702 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1607639953
transform 1 0 37610 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_434
timestamp 1607639953
transform 1 0 41014 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_422
timestamp 1607639953
transform 1 0 39910 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_459
timestamp 1607639953
transform 1 0 43314 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_446
timestamp 1607639953
transform 1 0 42118 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1607639953
transform 1 0 43222 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_483
timestamp 1607639953
transform 1 0 45522 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_471
timestamp 1607639953
transform 1 0 44418 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_495
timestamp 1607639953
transform 1 0 46626 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_520
timestamp 1607639953
transform 1 0 48926 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_507
timestamp 1607639953
transform 1 0 47730 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1607639953
transform 1 0 48834 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_544
timestamp 1607639953
transform 1 0 51134 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_532
timestamp 1607639953
transform 1 0 50030 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_568
timestamp 1607639953
transform 1 0 53342 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_556
timestamp 1607639953
transform 1 0 52238 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_593
timestamp 1607639953
transform 1 0 55642 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_581
timestamp 1607639953
transform 1 0 54538 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1607639953
transform 1 0 54446 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_605
timestamp 1607639953
transform 1 0 56746 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_617
timestamp 1607639953
transform 1 0 57850 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1607639953
transform -1 0 58862 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1607639953
transform 1 0 2466 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1607639953
transform 1 0 1362 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1607639953
transform 1 0 2466 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1607639953
transform 1 0 1362 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1607639953
transform 1 0 1086 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1607639953
transform 1 0 1086 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1607639953
transform 1 0 5134 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1607639953
transform 1 0 4030 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1607639953
transform 1 0 3570 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1607639953
transform 1 0 4674 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1607639953
transform 1 0 3570 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1607639953
transform 1 0 3938 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1607639953
transform 1 0 6238 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_62
timestamp 1607639953
transform 1 0 6790 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1607639953
transform 1 0 6514 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1607639953
transform 1 0 5778 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1607639953
transform 1 0 6698 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1607639953
transform 1 0 8446 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1607639953
transform 1 0 7342 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_84
timestamp 1607639953
transform 1 0 8814 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_72
timestamp 1607639953
transform 1 0 7710 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_68
timestamp 1607639953
transform 1 0 7342 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _097_
timestamp 1607639953
transform 1 0 7434 0 1 23392
box -38 -48 314 592
use OAI21X1  OAI21X1
timestamp 1608122862
transform 1 0 8078 0 1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1607639953
transform 1 0 10746 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1607639953
transform 1 0 9642 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_108
timestamp 1607639953
transform 1 0 11022 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_96
timestamp 1607639953
transform 1 0 9918 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1607639953
transform 1 0 9550 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1607639953
transform 1 0 12954 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_117
timestamp 1607639953
transform 1 0 11850 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_129
timestamp 1607639953
transform 1 0 12954 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_123
timestamp 1607639953
transform 1 0 12402 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_120
timestamp 1607639953
transform 1 0 12126 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1607639953
transform 1 0 12310 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _161_
timestamp 1607639953
transform 1 0 12678 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1607639953
transform 1 0 15254 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1607639953
transform 1 0 14058 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_153
timestamp 1607639953
transform 1 0 15162 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_141
timestamp 1607639953
transform 1 0 14058 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1607639953
transform 1 0 15162 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_166
timestamp 1607639953
transform 1 0 16358 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_165
timestamp 1607639953
transform 1 0 16266 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_190
timestamp 1607639953
transform 1 0 18566 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1607639953
transform 1 0 17462 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_187
timestamp 1607639953
transform 1 0 18290 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_177
timestamp 1607639953
transform 1 0 17370 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1607639953
transform 1 0 17922 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1607639953
transform 1 0 18014 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1607639953
transform 1 0 20866 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_202
timestamp 1607639953
transform 1 0 19670 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_218
timestamp 1607639953
transform 1 0 21142 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_206
timestamp 1607639953
transform 1 0 20038 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_199
timestamp 1607639953
transform 1 0 19394 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1607639953
transform 1 0 20774 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _207_
timestamp 1607639953
transform 1 0 19762 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1607639953
transform 1 0 23074 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1607639953
transform 1 0 21970 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_242
timestamp 1607639953
transform 1 0 23350 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_230
timestamp 1607639953
transform 1 0 22246 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_263
timestamp 1607639953
transform 1 0 25282 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_251
timestamp 1607639953
transform 1 0 24178 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_257
timestamp 1607639953
transform 1 0 24730 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1607639953
transform 1 0 23626 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1607639953
transform 1 0 23534 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_276
timestamp 1607639953
transform 1 0 26478 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1607639953
transform 1 0 26938 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_269
timestamp 1607639953
transform 1 0 25834 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1607639953
transform 1 0 26386 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_299
timestamp 1607639953
transform 1 0 28594 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_288
timestamp 1607639953
transform 1 0 27582 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_306
timestamp 1607639953
transform 1 0 29238 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1607639953
transform 1 0 28042 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1607639953
transform 1 0 29146 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _187_
timestamp 1607639953
transform 1 0 28318 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_323
timestamp 1607639953
transform 1 0 30802 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_311
timestamp 1607639953
transform 1 0 29698 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_330
timestamp 1607639953
transform 1 0 31446 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_318
timestamp 1607639953
transform 1 0 30342 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_349
timestamp 1607639953
transform 1 0 33194 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_337
timestamp 1607639953
transform 1 0 32090 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_335
timestamp 1607639953
transform 1 0 31906 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_342
timestamp 1607639953
transform 1 0 32550 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1607639953
transform 1 0 31998 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_373
timestamp 1607639953
transform 1 0 35402 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_361
timestamp 1607639953
transform 1 0 34298 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_367
timestamp 1607639953
transform 1 0 34850 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_354
timestamp 1607639953
transform 1 0 33654 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1607639953
transform 1 0 34758 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_385
timestamp 1607639953
transform 1 0 36506 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_391
timestamp 1607639953
transform 1 0 37058 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_379
timestamp 1607639953
transform 1 0 35954 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_410
timestamp 1607639953
transform 1 0 38806 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_398
timestamp 1607639953
transform 1 0 37702 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_415
timestamp 1607639953
transform 1 0 39266 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_403
timestamp 1607639953
transform 1 0 38162 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1607639953
transform 1 0 37610 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_434
timestamp 1607639953
transform 1 0 41014 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_422
timestamp 1607639953
transform 1 0 39910 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_440
timestamp 1607639953
transform 1 0 41566 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_428
timestamp 1607639953
transform 1 0 40462 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1607639953
transform 1 0 40370 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_459
timestamp 1607639953
transform 1 0 43314 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_446
timestamp 1607639953
transform 1 0 42118 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_452
timestamp 1607639953
transform 1 0 42670 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1607639953
transform 1 0 43222 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1607639953
transform 1 0 43406 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_475
timestamp 1607639953
transform 1 0 44786 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_463
timestamp 1607639953
transform 1 0 43682 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_476
timestamp 1607639953
transform 1 0 44878 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_464
timestamp 1607639953
transform 1 0 43774 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_499
timestamp 1607639953
transform 1 0 46994 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_487
timestamp 1607639953
transform 1 0 45890 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_501
timestamp 1607639953
transform 1 0 47178 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_489
timestamp 1607639953
transform 1 0 46074 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1607639953
transform 1 0 45982 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_520
timestamp 1607639953
transform 1 0 48926 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_511
timestamp 1607639953
transform 1 0 48098 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_525
timestamp 1607639953
transform 1 0 49386 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_513
timestamp 1607639953
transform 1 0 48282 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1607639953
transform 1 0 48834 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_544
timestamp 1607639953
transform 1 0 51134 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_532
timestamp 1607639953
transform 1 0 50030 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_550
timestamp 1607639953
transform 1 0 51686 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_537
timestamp 1607639953
transform 1 0 50490 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1607639953
transform 1 0 51594 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_568
timestamp 1607639953
transform 1 0 53342 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_556
timestamp 1607639953
transform 1 0 52238 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_562
timestamp 1607639953
transform 1 0 52790 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_593
timestamp 1607639953
transform 1 0 55642 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_581
timestamp 1607639953
transform 1 0 54538 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_586
timestamp 1607639953
transform 1 0 54998 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_574
timestamp 1607639953
transform 1 0 53894 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1607639953
transform 1 0 54446 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_605
timestamp 1607639953
transform 1 0 56746 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_611
timestamp 1607639953
transform 1 0 57298 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_598
timestamp 1607639953
transform 1 0 56102 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1607639953
transform 1 0 57206 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_617
timestamp 1607639953
transform 1 0 57850 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_623
timestamp 1607639953
transform 1 0 58402 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1607639953
transform -1 0 58862 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1607639953
transform -1 0 58862 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_16
timestamp 1607639953
transform 1 0 2558 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1607639953
transform 1 0 2098 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_3
timestamp 1607639953
transform 1 0 1362 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1607639953
transform 1 0 1086 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _103_
timestamp 1607639953
transform 1 0 2282 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_40
timestamp 1607639953
transform 1 0 4766 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_28
timestamp 1607639953
transform 1 0 3662 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1607639953
transform 1 0 6790 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_60
timestamp 1607639953
transform 1 0 6606 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_52
timestamp 1607639953
transform 1 0 5870 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1607639953
transform 1 0 6698 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1607639953
transform 1 0 8998 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_74
timestamp 1607639953
transform 1 0 7894 0 1 24480
box -38 -48 222 592
use OAI22X1  OAI22X1
timestamp 1608122862
transform 1 0 8078 0 1 24480
box 0 -48 920 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1607639953
transform 1 0 11206 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1607639953
transform 1 0 10102 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1607639953
transform 1 0 12402 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1607639953
transform 1 0 12310 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_147
timestamp 1607639953
transform 1 0 14610 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1607639953
transform 1 0 13506 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_171
timestamp 1607639953
transform 1 0 16818 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_159
timestamp 1607639953
transform 1 0 15714 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1607639953
transform 1 0 19118 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1607639953
transform 1 0 18014 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1607639953
transform 1 0 17922 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1607639953
transform 1 0 21326 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1607639953
transform 1 0 20222 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1607639953
transform 1 0 22430 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1607639953
transform 1 0 24730 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1607639953
transform 1 0 23626 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1607639953
transform 1 0 23534 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1607639953
transform 1 0 26938 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_269
timestamp 1607639953
transform 1 0 25834 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_306
timestamp 1607639953
transform 1 0 29238 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1607639953
transform 1 0 28042 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1607639953
transform 1 0 29146 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_330
timestamp 1607639953
transform 1 0 31446 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_318
timestamp 1607639953
transform 1 0 30342 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_342
timestamp 1607639953
transform 1 0 32550 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_367
timestamp 1607639953
transform 1 0 34850 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_354
timestamp 1607639953
transform 1 0 33654 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1607639953
transform 1 0 34758 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_391
timestamp 1607639953
transform 1 0 37058 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_379
timestamp 1607639953
transform 1 0 35954 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_415
timestamp 1607639953
transform 1 0 39266 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_403
timestamp 1607639953
transform 1 0 38162 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_440
timestamp 1607639953
transform 1 0 41566 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_428
timestamp 1607639953
transform 1 0 40462 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1607639953
transform 1 0 40370 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_452
timestamp 1607639953
transform 1 0 42670 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_476
timestamp 1607639953
transform 1 0 44878 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_464
timestamp 1607639953
transform 1 0 43774 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_501
timestamp 1607639953
transform 1 0 47178 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_489
timestamp 1607639953
transform 1 0 46074 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1607639953
transform 1 0 45982 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_525
timestamp 1607639953
transform 1 0 49386 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_513
timestamp 1607639953
transform 1 0 48282 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_550
timestamp 1607639953
transform 1 0 51686 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_537
timestamp 1607639953
transform 1 0 50490 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1607639953
transform 1 0 51594 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_562
timestamp 1607639953
transform 1 0 52790 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_586
timestamp 1607639953
transform 1 0 54998 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_574
timestamp 1607639953
transform 1 0 53894 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_611
timestamp 1607639953
transform 1 0 57298 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_598
timestamp 1607639953
transform 1 0 56102 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1607639953
transform 1 0 57206 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_623
timestamp 1607639953
transform 1 0 58402 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1607639953
transform -1 0 58862 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1607639953
transform 1 0 2466 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1607639953
transform 1 0 1362 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1607639953
transform 1 0 1086 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1607639953
transform 1 0 5134 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1607639953
transform 1 0 4030 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1607639953
transform 1 0 3570 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1607639953
transform 1 0 3938 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_56
timestamp 1607639953
transform 1 0 6238 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_80
timestamp 1607639953
transform 1 0 8446 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_68
timestamp 1607639953
transform 1 0 7342 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_105
timestamp 1607639953
transform 1 0 10746 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_93
timestamp 1607639953
transform 1 0 9642 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1607639953
transform 1 0 9550 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_129
timestamp 1607639953
transform 1 0 12954 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_117
timestamp 1607639953
transform 1 0 11850 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_154
timestamp 1607639953
transform 1 0 15254 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1607639953
transform 1 0 14058 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1607639953
transform 1 0 15162 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_166
timestamp 1607639953
transform 1 0 16358 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_190
timestamp 1607639953
transform 1 0 18566 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_178
timestamp 1607639953
transform 1 0 17462 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_215
timestamp 1607639953
transform 1 0 20866 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_202
timestamp 1607639953
transform 1 0 19670 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1607639953
transform 1 0 20774 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_239
timestamp 1607639953
transform 1 0 23074 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_227
timestamp 1607639953
transform 1 0 21970 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_263
timestamp 1607639953
transform 1 0 25282 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_251
timestamp 1607639953
transform 1 0 24178 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_276
timestamp 1607639953
transform 1 0 26478 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1607639953
transform 1 0 26386 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_300
timestamp 1607639953
transform 1 0 28686 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_288
timestamp 1607639953
transform 1 0 27582 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_324
timestamp 1607639953
transform 1 0 30894 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_312
timestamp 1607639953
transform 1 0 29790 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_349
timestamp 1607639953
transform 1 0 33194 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_337
timestamp 1607639953
transform 1 0 32090 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1607639953
transform 1 0 31998 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_373
timestamp 1607639953
transform 1 0 35402 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_361
timestamp 1607639953
transform 1 0 34298 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_385
timestamp 1607639953
transform 1 0 36506 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_410
timestamp 1607639953
transform 1 0 38806 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_398
timestamp 1607639953
transform 1 0 37702 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1607639953
transform 1 0 37610 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_434
timestamp 1607639953
transform 1 0 41014 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_422
timestamp 1607639953
transform 1 0 39910 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_459
timestamp 1607639953
transform 1 0 43314 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_446
timestamp 1607639953
transform 1 0 42118 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1607639953
transform 1 0 43222 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_483
timestamp 1607639953
transform 1 0 45522 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_471
timestamp 1607639953
transform 1 0 44418 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_495
timestamp 1607639953
transform 1 0 46626 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_520
timestamp 1607639953
transform 1 0 48926 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_507
timestamp 1607639953
transform 1 0 47730 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1607639953
transform 1 0 48834 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_544
timestamp 1607639953
transform 1 0 51134 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_532
timestamp 1607639953
transform 1 0 50030 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _093_
timestamp 1607639953
transform 1 0 51502 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_563
timestamp 1607639953
transform 1 0 52882 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_551
timestamp 1607639953
transform 1 0 51778 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_593
timestamp 1607639953
transform 1 0 55642 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_581
timestamp 1607639953
transform 1 0 54538 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_579
timestamp 1607639953
transform 1 0 54354 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_575
timestamp 1607639953
transform 1 0 53986 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1607639953
transform 1 0 54446 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_605
timestamp 1607639953
transform 1 0 56746 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_617
timestamp 1607639953
transform 1 0 57850 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1607639953
transform -1 0 58862 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1607639953
transform 1 0 2466 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1607639953
transform 1 0 1362 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1607639953
transform 1 0 1086 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1607639953
transform 1 0 4674 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1607639953
transform 1 0 3570 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_62
timestamp 1607639953
transform 1 0 6790 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_59
timestamp 1607639953
transform 1 0 6514 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_51
timestamp 1607639953
transform 1 0 5778 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1607639953
transform 1 0 6698 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_84
timestamp 1607639953
transform 1 0 8814 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_74
timestamp 1607639953
transform 1 0 7894 0 1 25568
box -38 -48 222 592
use OR2X1  OR2X1
timestamp 1608122862
transform 1 0 8078 0 1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_43_100
timestamp 1607639953
transform 1 0 10286 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_96
timestamp 1607639953
transform 1 0 9918 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _163_
timestamp 1607639953
transform 1 0 10010 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_131
timestamp 1607639953
transform 1 0 13138 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_123
timestamp 1607639953
transform 1 0 12402 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_120
timestamp 1607639953
transform 1 0 12126 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_112
timestamp 1607639953
transform 1 0 11390 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1607639953
transform 1 0 12310 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1607639953
transform 1 0 14794 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1607639953
transform 1 0 13690 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1607639953
transform 1 0 13414 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_173
timestamp 1607639953
transform 1 0 17002 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_161
timestamp 1607639953
transform 1 0 15898 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_196
timestamp 1607639953
transform 1 0 19118 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_184
timestamp 1607639953
transform 1 0 18014 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_181
timestamp 1607639953
transform 1 0 17738 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1607639953
transform 1 0 17922 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_220
timestamp 1607639953
transform 1 0 21326 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_208
timestamp 1607639953
transform 1 0 20222 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_232
timestamp 1607639953
transform 1 0 22430 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_257
timestamp 1607639953
transform 1 0 24730 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_245
timestamp 1607639953
transform 1 0 23626 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1607639953
transform 1 0 23534 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1607639953
transform 1 0 26938 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_269
timestamp 1607639953
transform 1 0 25834 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_306
timestamp 1607639953
transform 1 0 29238 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1607639953
transform 1 0 28042 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1607639953
transform 1 0 29146 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_330
timestamp 1607639953
transform 1 0 31446 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_318
timestamp 1607639953
transform 1 0 30342 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_342
timestamp 1607639953
transform 1 0 32550 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_367
timestamp 1607639953
transform 1 0 34850 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_354
timestamp 1607639953
transform 1 0 33654 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1607639953
transform 1 0 34758 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_391
timestamp 1607639953
transform 1 0 37058 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_379
timestamp 1607639953
transform 1 0 35954 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_415
timestamp 1607639953
transform 1 0 39266 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_403
timestamp 1607639953
transform 1 0 38162 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_440
timestamp 1607639953
transform 1 0 41566 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_428
timestamp 1607639953
transform 1 0 40462 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1607639953
transform 1 0 40370 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_460
timestamp 1607639953
transform 1 0 43406 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_448
timestamp 1607639953
transform 1 0 42302 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_444
timestamp 1607639953
transform 1 0 41934 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _072_
timestamp 1607639953
transform 1 0 42026 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_484
timestamp 1607639953
transform 1 0 45614 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_472
timestamp 1607639953
transform 1 0 44510 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_501
timestamp 1607639953
transform 1 0 47178 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_489
timestamp 1607639953
transform 1 0 46074 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1607639953
transform 1 0 45982 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_525
timestamp 1607639953
transform 1 0 49386 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_513
timestamp 1607639953
transform 1 0 48282 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_550
timestamp 1607639953
transform 1 0 51686 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_537
timestamp 1607639953
transform 1 0 50490 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1607639953
transform 1 0 51594 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_562
timestamp 1607639953
transform 1 0 52790 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_586
timestamp 1607639953
transform 1 0 54998 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_574
timestamp 1607639953
transform 1 0 53894 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_611
timestamp 1607639953
transform 1 0 57298 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_598
timestamp 1607639953
transform 1 0 56102 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1607639953
transform 1 0 57206 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_623
timestamp 1607639953
transform 1 0 58402 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1607639953
transform -1 0 58862 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1607639953
transform 1 0 2466 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1607639953
transform 1 0 1362 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1607639953
transform 1 0 1086 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_44
timestamp 1607639953
transform 1 0 5134 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_32
timestamp 1607639953
transform 1 0 4030 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1607639953
transform 1 0 3570 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1607639953
transform 1 0 3938 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_56
timestamp 1607639953
transform 1 0 6238 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_80
timestamp 1607639953
transform 1 0 8446 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_68
timestamp 1607639953
transform 1 0 7342 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_105
timestamp 1607639953
transform 1 0 10746 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_93
timestamp 1607639953
transform 1 0 9642 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1607639953
transform 1 0 9550 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_129
timestamp 1607639953
transform 1 0 12954 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_117
timestamp 1607639953
transform 1 0 11850 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_154
timestamp 1607639953
transform 1 0 15254 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1607639953
transform 1 0 14058 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1607639953
transform 1 0 15162 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_166
timestamp 1607639953
transform 1 0 16358 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_190
timestamp 1607639953
transform 1 0 18566 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_178
timestamp 1607639953
transform 1 0 17462 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_215
timestamp 1607639953
transform 1 0 20866 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_202
timestamp 1607639953
transform 1 0 19670 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1607639953
transform 1 0 20774 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_239
timestamp 1607639953
transform 1 0 23074 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_227
timestamp 1607639953
transform 1 0 21970 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_261
timestamp 1607639953
transform 1 0 25098 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_257
timestamp 1607639953
transform 1 0 24730 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_251
timestamp 1607639953
transform 1 0 24178 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _137_
timestamp 1607639953
transform 1 0 24822 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_276
timestamp 1607639953
transform 1 0 26478 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_273
timestamp 1607639953
transform 1 0 26202 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1607639953
transform 1 0 26386 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_308
timestamp 1607639953
transform 1 0 29422 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_304
timestamp 1607639953
transform 1 0 29054 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_300
timestamp 1607639953
transform 1 0 28686 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_288
timestamp 1607639953
transform 1 0 27582 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _019_
timestamp 1607639953
transform 1 0 29146 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_320
timestamp 1607639953
transform 1 0 30526 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_349
timestamp 1607639953
transform 1 0 33194 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_337
timestamp 1607639953
transform 1 0 32090 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_332
timestamp 1607639953
transform 1 0 31630 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1607639953
transform 1 0 31998 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_372
timestamp 1607639953
transform 1 0 35310 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_360
timestamp 1607639953
transform 1 0 34206 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _095_
timestamp 1607639953
transform 1 0 33930 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_396
timestamp 1607639953
transform 1 0 37518 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_384
timestamp 1607639953
transform 1 0 36414 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_410
timestamp 1607639953
transform 1 0 38806 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_398
timestamp 1607639953
transform 1 0 37702 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1607639953
transform 1 0 37610 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_434
timestamp 1607639953
transform 1 0 41014 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_422
timestamp 1607639953
transform 1 0 39910 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_462
timestamp 1607639953
transform 1 0 43590 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_446
timestamp 1607639953
transform 1 0 42118 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1607639953
transform 1 0 43222 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _188_
timestamp 1607639953
transform 1 0 43314 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_474
timestamp 1607639953
transform 1 0 44694 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_498
timestamp 1607639953
transform 1 0 46902 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_486
timestamp 1607639953
transform 1 0 45798 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_523
timestamp 1607639953
transform 1 0 49202 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_518
timestamp 1607639953
transform 1 0 48742 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_510
timestamp 1607639953
transform 1 0 48006 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1607639953
transform 1 0 48834 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _096_
timestamp 1607639953
transform 1 0 48926 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_547
timestamp 1607639953
transform 1 0 51410 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_535
timestamp 1607639953
transform 1 0 50306 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_571
timestamp 1607639953
transform 1 0 53618 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_559
timestamp 1607639953
transform 1 0 52514 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_593
timestamp 1607639953
transform 1 0 55642 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_581
timestamp 1607639953
transform 1 0 54538 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_579
timestamp 1607639953
transform 1 0 54354 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1607639953
transform 1 0 54446 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_605
timestamp 1607639953
transform 1 0 56746 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_617
timestamp 1607639953
transform 1 0 57850 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1607639953
transform -1 0 58862 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1607639953
transform 1 0 2466 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1607639953
transform 1 0 1362 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1607639953
transform 1 0 1086 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1607639953
transform 1 0 4674 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1607639953
transform 1 0 3570 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_62
timestamp 1607639953
transform 1 0 6790 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_59
timestamp 1607639953
transform 1 0 6514 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_51
timestamp 1607639953
transform 1 0 5778 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1607639953
transform 1 0 6698 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_84
timestamp 1607639953
transform 1 0 8814 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_74
timestamp 1607639953
transform 1 0 7894 0 1 26656
box -38 -48 222 592
use OR2X2  OR2X2
timestamp 1608122862
transform 1 0 8078 0 1 26656
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_45_108
timestamp 1607639953
transform 1 0 11022 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_96
timestamp 1607639953
transform 1 0 9918 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_123
timestamp 1607639953
transform 1 0 12402 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_120
timestamp 1607639953
transform 1 0 12126 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1607639953
transform 1 0 12310 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_147
timestamp 1607639953
transform 1 0 14610 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_135
timestamp 1607639953
transform 1 0 13506 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_171
timestamp 1607639953
transform 1 0 16818 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_159
timestamp 1607639953
transform 1 0 15714 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_196
timestamp 1607639953
transform 1 0 19118 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_184
timestamp 1607639953
transform 1 0 18014 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1607639953
transform 1 0 17922 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1607639953
transform 1 0 21326 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_208
timestamp 1607639953
transform 1 0 20222 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_239
timestamp 1607639953
transform 1 0 23074 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_227
timestamp 1607639953
transform 1 0 21970 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _009_
timestamp 1607639953
transform 1 0 21694 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_257
timestamp 1607639953
transform 1 0 24730 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_245
timestamp 1607639953
transform 1 0 23626 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_243
timestamp 1607639953
transform 1 0 23442 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1607639953
transform 1 0 23534 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1607639953
transform 1 0 26938 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_269
timestamp 1607639953
transform 1 0 25834 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_306
timestamp 1607639953
transform 1 0 29238 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1607639953
transform 1 0 28042 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1607639953
transform 1 0 29146 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_330
timestamp 1607639953
transform 1 0 31446 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_318
timestamp 1607639953
transform 1 0 30342 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_342
timestamp 1607639953
transform 1 0 32550 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_367
timestamp 1607639953
transform 1 0 34850 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_354
timestamp 1607639953
transform 1 0 33654 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1607639953
transform 1 0 34758 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_391
timestamp 1607639953
transform 1 0 37058 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_379
timestamp 1607639953
transform 1 0 35954 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_414
timestamp 1607639953
transform 1 0 39174 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_402
timestamp 1607639953
transform 1 0 38070 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _081_
timestamp 1607639953
transform 1 0 37794 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_440
timestamp 1607639953
transform 1 0 41566 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_428
timestamp 1607639953
transform 1 0 40462 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_426
timestamp 1607639953
transform 1 0 40278 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1607639953
transform 1 0 40370 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_452
timestamp 1607639953
transform 1 0 42670 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_476
timestamp 1607639953
transform 1 0 44878 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_464
timestamp 1607639953
transform 1 0 43774 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_501
timestamp 1607639953
transform 1 0 47178 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_489
timestamp 1607639953
transform 1 0 46074 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1607639953
transform 1 0 45982 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_525
timestamp 1607639953
transform 1 0 49386 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_513
timestamp 1607639953
transform 1 0 48282 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_550
timestamp 1607639953
transform 1 0 51686 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_537
timestamp 1607639953
transform 1 0 50490 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1607639953
transform 1 0 51594 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_562
timestamp 1607639953
transform 1 0 52790 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_586
timestamp 1607639953
transform 1 0 54998 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_574
timestamp 1607639953
transform 1 0 53894 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_611
timestamp 1607639953
transform 1 0 57298 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_598
timestamp 1607639953
transform 1 0 56102 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1607639953
transform 1 0 57206 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_623
timestamp 1607639953
transform 1 0 58402 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1607639953
transform -1 0 58862 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1607639953
transform 1 0 2466 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1607639953
transform 1 0 1362 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1607639953
transform 1 0 2466 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1607639953
transform 1 0 1362 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1607639953
transform 1 0 1086 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1607639953
transform 1 0 1086 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1607639953
transform 1 0 4674 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1607639953
transform 1 0 3570 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_44
timestamp 1607639953
transform 1 0 5134 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_32
timestamp 1607639953
transform 1 0 4030 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_27
timestamp 1607639953
transform 1 0 3570 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1607639953
transform 1 0 3938 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_62
timestamp 1607639953
transform 1 0 6790 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_59
timestamp 1607639953
transform 1 0 6514 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_51
timestamp 1607639953
transform 1 0 5778 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_56
timestamp 1607639953
transform 1 0 6238 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1607639953
transform 1 0 6698 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_84
timestamp 1607639953
transform 1 0 8814 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_74
timestamp 1607639953
transform 1 0 7894 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_80
timestamp 1607639953
transform 1 0 8446 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_68
timestamp 1607639953
transform 1 0 7342 0 -1 27744
box -38 -48 1142 592
use TBUFX1  TBUFX1
timestamp 1608122862
transform 1 0 8078 0 1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_47_108
timestamp 1607639953
transform 1 0 11022 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_96
timestamp 1607639953
transform 1 0 9918 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_105
timestamp 1607639953
transform 1 0 10746 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_93
timestamp 1607639953
transform 1 0 9642 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1607639953
transform 1 0 9550 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_123
timestamp 1607639953
transform 1 0 12402 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_120
timestamp 1607639953
transform 1 0 12126 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_129
timestamp 1607639953
transform 1 0 12954 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_117
timestamp 1607639953
transform 1 0 11850 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1607639953
transform 1 0 12310 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_147
timestamp 1607639953
transform 1 0 14610 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_135
timestamp 1607639953
transform 1 0 13506 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_154
timestamp 1607639953
transform 1 0 15254 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1607639953
transform 1 0 14058 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1607639953
transform 1 0 15162 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_171
timestamp 1607639953
transform 1 0 16818 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_159
timestamp 1607639953
transform 1 0 15714 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_166
timestamp 1607639953
transform 1 0 16358 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_196
timestamp 1607639953
transform 1 0 19118 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_184
timestamp 1607639953
transform 1 0 18014 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_190
timestamp 1607639953
transform 1 0 18566 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_178
timestamp 1607639953
transform 1 0 17462 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1607639953
transform 1 0 17922 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_220
timestamp 1607639953
transform 1 0 21326 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_208
timestamp 1607639953
transform 1 0 20222 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_215
timestamp 1607639953
transform 1 0 20866 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_202
timestamp 1607639953
transform 1 0 19670 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1607639953
transform 1 0 20774 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_232
timestamp 1607639953
transform 1 0 22430 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_239
timestamp 1607639953
transform 1 0 23074 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_227
timestamp 1607639953
transform 1 0 21970 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_257
timestamp 1607639953
transform 1 0 24730 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_245
timestamp 1607639953
transform 1 0 23626 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_263
timestamp 1607639953
transform 1 0 25282 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_251
timestamp 1607639953
transform 1 0 24178 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1607639953
transform 1 0 23534 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1607639953
transform 1 0 26938 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_269
timestamp 1607639953
transform 1 0 25834 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_276
timestamp 1607639953
transform 1 0 26478 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1607639953
transform 1 0 26386 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_306
timestamp 1607639953
transform 1 0 29238 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1607639953
transform 1 0 28042 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_300
timestamp 1607639953
transform 1 0 28686 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_288
timestamp 1607639953
transform 1 0 27582 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1607639953
transform 1 0 29146 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_330
timestamp 1607639953
transform 1 0 31446 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_318
timestamp 1607639953
transform 1 0 30342 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_324
timestamp 1607639953
transform 1 0 30894 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_312
timestamp 1607639953
transform 1 0 29790 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_342
timestamp 1607639953
transform 1 0 32550 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_349
timestamp 1607639953
transform 1 0 33194 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_337
timestamp 1607639953
transform 1 0 32090 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1607639953
transform 1 0 31998 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_367
timestamp 1607639953
transform 1 0 34850 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_354
timestamp 1607639953
transform 1 0 33654 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_373
timestamp 1607639953
transform 1 0 35402 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_361
timestamp 1607639953
transform 1 0 34298 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1607639953
transform 1 0 34758 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_391
timestamp 1607639953
transform 1 0 37058 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_379
timestamp 1607639953
transform 1 0 35954 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_385
timestamp 1607639953
transform 1 0 36506 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_412
timestamp 1607639953
transform 1 0 38990 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_400
timestamp 1607639953
transform 1 0 37886 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_410
timestamp 1607639953
transform 1 0 38806 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_398
timestamp 1607639953
transform 1 0 37702 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1607639953
transform 1 0 37610 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _142_
timestamp 1607639953
transform 1 0 37610 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_440
timestamp 1607639953
transform 1 0 41566 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_428
timestamp 1607639953
transform 1 0 40462 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_424
timestamp 1607639953
transform 1 0 40094 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_434
timestamp 1607639953
transform 1 0 41014 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_422
timestamp 1607639953
transform 1 0 39910 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1607639953
transform 1 0 40370 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_452
timestamp 1607639953
transform 1 0 42670 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_459
timestamp 1607639953
transform 1 0 43314 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_446
timestamp 1607639953
transform 1 0 42118 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1607639953
transform 1 0 43222 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_476
timestamp 1607639953
transform 1 0 44878 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_464
timestamp 1607639953
transform 1 0 43774 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_483
timestamp 1607639953
transform 1 0 45522 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_471
timestamp 1607639953
transform 1 0 44418 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_501
timestamp 1607639953
transform 1 0 47178 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_489
timestamp 1607639953
transform 1 0 46074 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_495
timestamp 1607639953
transform 1 0 46626 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1607639953
transform 1 0 45982 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_525
timestamp 1607639953
transform 1 0 49386 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_513
timestamp 1607639953
transform 1 0 48282 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_520
timestamp 1607639953
transform 1 0 48926 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_507
timestamp 1607639953
transform 1 0 47730 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1607639953
transform 1 0 48834 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_550
timestamp 1607639953
transform 1 0 51686 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_537
timestamp 1607639953
transform 1 0 50490 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_544
timestamp 1607639953
transform 1 0 51134 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_532
timestamp 1607639953
transform 1 0 50030 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1607639953
transform 1 0 51594 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_562
timestamp 1607639953
transform 1 0 52790 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_568
timestamp 1607639953
transform 1 0 53342 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_556
timestamp 1607639953
transform 1 0 52238 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_586
timestamp 1607639953
transform 1 0 54998 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_574
timestamp 1607639953
transform 1 0 53894 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_593
timestamp 1607639953
transform 1 0 55642 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_581
timestamp 1607639953
transform 1 0 54538 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1607639953
transform 1 0 54446 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_611
timestamp 1607639953
transform 1 0 57298 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_598
timestamp 1607639953
transform 1 0 56102 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_605
timestamp 1607639953
transform 1 0 56746 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1607639953
transform 1 0 57206 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_623
timestamp 1607639953
transform 1 0 58402 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_617
timestamp 1607639953
transform 1 0 57850 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1607639953
transform -1 0 58862 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1607639953
transform -1 0 58862 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1607639953
transform 1 0 2466 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1607639953
transform 1 0 1362 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1607639953
transform 1 0 1086 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_44
timestamp 1607639953
transform 1 0 5134 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_32
timestamp 1607639953
transform 1 0 4030 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_27
timestamp 1607639953
transform 1 0 3570 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1607639953
transform 1 0 3938 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_56
timestamp 1607639953
transform 1 0 6238 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_80
timestamp 1607639953
transform 1 0 8446 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_68
timestamp 1607639953
transform 1 0 7342 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_105
timestamp 1607639953
transform 1 0 10746 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_93
timestamp 1607639953
transform 1 0 9642 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1607639953
transform 1 0 9550 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_129
timestamp 1607639953
transform 1 0 12954 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_117
timestamp 1607639953
transform 1 0 11850 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_154
timestamp 1607639953
transform 1 0 15254 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1607639953
transform 1 0 14058 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1607639953
transform 1 0 15162 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_166
timestamp 1607639953
transform 1 0 16358 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_190
timestamp 1607639953
transform 1 0 18566 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_178
timestamp 1607639953
transform 1 0 17462 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_215
timestamp 1607639953
transform 1 0 20866 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_202
timestamp 1607639953
transform 1 0 19670 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1607639953
transform 1 0 20774 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_239
timestamp 1607639953
transform 1 0 23074 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_227
timestamp 1607639953
transform 1 0 21970 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_263
timestamp 1607639953
transform 1 0 25282 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_251
timestamp 1607639953
transform 1 0 24178 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_276
timestamp 1607639953
transform 1 0 26478 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_271
timestamp 1607639953
transform 1 0 26018 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_267
timestamp 1607639953
transform 1 0 25650 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1607639953
transform 1 0 26386 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _206_
timestamp 1607639953
transform 1 0 25742 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_303
timestamp 1607639953
transform 1 0 28962 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_291
timestamp 1607639953
transform 1 0 27858 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _006_
timestamp 1607639953
transform 1 0 27582 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_327
timestamp 1607639953
transform 1 0 31170 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_315
timestamp 1607639953
transform 1 0 30066 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_349
timestamp 1607639953
transform 1 0 33194 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_337
timestamp 1607639953
transform 1 0 32090 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_335
timestamp 1607639953
transform 1 0 31906 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1607639953
transform 1 0 31998 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_367
timestamp 1607639953
transform 1 0 34850 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_361
timestamp 1607639953
transform 1 0 34298 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _204_
timestamp 1607639953
transform 1 0 34574 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_391
timestamp 1607639953
transform 1 0 37058 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_379
timestamp 1607639953
transform 1 0 35954 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_410
timestamp 1607639953
transform 1 0 38806 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_398
timestamp 1607639953
transform 1 0 37702 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1607639953
transform 1 0 37610 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_434
timestamp 1607639953
transform 1 0 41014 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_422
timestamp 1607639953
transform 1 0 39910 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_459
timestamp 1607639953
transform 1 0 43314 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_446
timestamp 1607639953
transform 1 0 42118 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1607639953
transform 1 0 43222 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_483
timestamp 1607639953
transform 1 0 45522 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_471
timestamp 1607639953
transform 1 0 44418 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_495
timestamp 1607639953
transform 1 0 46626 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_520
timestamp 1607639953
transform 1 0 48926 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_507
timestamp 1607639953
transform 1 0 47730 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1607639953
transform 1 0 48834 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_544
timestamp 1607639953
transform 1 0 51134 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_532
timestamp 1607639953
transform 1 0 50030 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_568
timestamp 1607639953
transform 1 0 53342 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_556
timestamp 1607639953
transform 1 0 52238 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_593
timestamp 1607639953
transform 1 0 55642 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_581
timestamp 1607639953
transform 1 0 54538 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1607639953
transform 1 0 54446 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_605
timestamp 1607639953
transform 1 0 56746 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_617
timestamp 1607639953
transform 1 0 57850 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1607639953
transform -1 0 58862 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_15
timestamp 1607639953
transform 1 0 2466 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1607639953
transform 1 0 1362 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1607639953
transform 1 0 1086 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_40
timestamp 1607639953
transform 1 0 4766 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_28
timestamp 1607639953
transform 1 0 3662 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_23
timestamp 1607639953
transform 1 0 3202 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _098_
timestamp 1607639953
transform 1 0 3386 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_62
timestamp 1607639953
transform 1 0 6790 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_60
timestamp 1607639953
transform 1 0 6606 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_52
timestamp 1607639953
transform 1 0 5870 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1607639953
transform 1 0 6698 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_88
timestamp 1607639953
transform 1 0 9182 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_74
timestamp 1607639953
transform 1 0 7894 0 1 28832
box -38 -48 222 592
use TBUFX2  TBUFX2
timestamp 1608122862
transform 1 0 8078 0 1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_49_100
timestamp 1607639953
transform 1 0 10286 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_123
timestamp 1607639953
transform 1 0 12402 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_120
timestamp 1607639953
transform 1 0 12126 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_112
timestamp 1607639953
transform 1 0 11390 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1607639953
transform 1 0 12310 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_147
timestamp 1607639953
transform 1 0 14610 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_135
timestamp 1607639953
transform 1 0 13506 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_171
timestamp 1607639953
transform 1 0 16818 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_159
timestamp 1607639953
transform 1 0 15714 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_196
timestamp 1607639953
transform 1 0 19118 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_184
timestamp 1607639953
transform 1 0 18014 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1607639953
transform 1 0 17922 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_220
timestamp 1607639953
transform 1 0 21326 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_208
timestamp 1607639953
transform 1 0 20222 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_232
timestamp 1607639953
transform 1 0 22430 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_257
timestamp 1607639953
transform 1 0 24730 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_245
timestamp 1607639953
transform 1 0 23626 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1607639953
transform 1 0 23534 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1607639953
transform 1 0 26938 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_269
timestamp 1607639953
transform 1 0 25834 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_306
timestamp 1607639953
transform 1 0 29238 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1607639953
transform 1 0 28042 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1607639953
transform 1 0 29146 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_319
timestamp 1607639953
transform 1 0 30434 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_314
timestamp 1607639953
transform 1 0 29974 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _201_
timestamp 1607639953
transform 1 0 30158 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_343
timestamp 1607639953
transform 1 0 32642 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_331
timestamp 1607639953
transform 1 0 31538 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_367
timestamp 1607639953
transform 1 0 34850 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_363
timestamp 1607639953
transform 1 0 34482 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_355
timestamp 1607639953
transform 1 0 33746 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1607639953
transform 1 0 34758 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_391
timestamp 1607639953
transform 1 0 37058 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_379
timestamp 1607639953
transform 1 0 35954 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_415
timestamp 1607639953
transform 1 0 39266 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_403
timestamp 1607639953
transform 1 0 38162 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_440
timestamp 1607639953
transform 1 0 41566 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_428
timestamp 1607639953
transform 1 0 40462 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1607639953
transform 1 0 40370 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_452
timestamp 1607639953
transform 1 0 42670 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_476
timestamp 1607639953
transform 1 0 44878 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_464
timestamp 1607639953
transform 1 0 43774 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_501
timestamp 1607639953
transform 1 0 47178 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_489
timestamp 1607639953
transform 1 0 46074 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1607639953
transform 1 0 45982 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_525
timestamp 1607639953
transform 1 0 49386 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_513
timestamp 1607639953
transform 1 0 48282 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_550
timestamp 1607639953
transform 1 0 51686 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_537
timestamp 1607639953
transform 1 0 50490 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1607639953
transform 1 0 51594 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_562
timestamp 1607639953
transform 1 0 52790 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_586
timestamp 1607639953
transform 1 0 54998 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_574
timestamp 1607639953
transform 1 0 53894 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_611
timestamp 1607639953
transform 1 0 57298 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_598
timestamp 1607639953
transform 1 0 56102 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1607639953
transform 1 0 57206 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_623
timestamp 1607639953
transform 1 0 58402 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1607639953
transform -1 0 58862 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1607639953
transform 1 0 2466 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1607639953
transform 1 0 1362 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1607639953
transform 1 0 1086 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_44
timestamp 1607639953
transform 1 0 5134 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_32
timestamp 1607639953
transform 1 0 4030 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_27
timestamp 1607639953
transform 1 0 3570 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1607639953
transform 1 0 3938 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_56
timestamp 1607639953
transform 1 0 6238 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_80
timestamp 1607639953
transform 1 0 8446 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_68
timestamp 1607639953
transform 1 0 7342 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_105
timestamp 1607639953
transform 1 0 10746 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_93
timestamp 1607639953
transform 1 0 9642 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1607639953
transform 1 0 9550 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_129
timestamp 1607639953
transform 1 0 12954 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_117
timestamp 1607639953
transform 1 0 11850 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_154
timestamp 1607639953
transform 1 0 15254 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1607639953
transform 1 0 14058 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1607639953
transform 1 0 15162 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_171
timestamp 1607639953
transform 1 0 16818 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_159
timestamp 1607639953
transform 1 0 15714 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _120_
timestamp 1607639953
transform 1 0 15438 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_195
timestamp 1607639953
transform 1 0 19026 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_183
timestamp 1607639953
transform 1 0 17922 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_215
timestamp 1607639953
transform 1 0 20866 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_213
timestamp 1607639953
transform 1 0 20682 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_207
timestamp 1607639953
transform 1 0 20130 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1607639953
transform 1 0 20774 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_239
timestamp 1607639953
transform 1 0 23074 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_227
timestamp 1607639953
transform 1 0 21970 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_263
timestamp 1607639953
transform 1 0 25282 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_251
timestamp 1607639953
transform 1 0 24178 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_276
timestamp 1607639953
transform 1 0 26478 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1607639953
transform 1 0 26386 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_300
timestamp 1607639953
transform 1 0 28686 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_288
timestamp 1607639953
transform 1 0 27582 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_324
timestamp 1607639953
transform 1 0 30894 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_312
timestamp 1607639953
transform 1 0 29790 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_349
timestamp 1607639953
transform 1 0 33194 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_337
timestamp 1607639953
transform 1 0 32090 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1607639953
transform 1 0 31998 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_373
timestamp 1607639953
transform 1 0 35402 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_361
timestamp 1607639953
transform 1 0 34298 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_385
timestamp 1607639953
transform 1 0 36506 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_410
timestamp 1607639953
transform 1 0 38806 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_398
timestamp 1607639953
transform 1 0 37702 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1607639953
transform 1 0 37610 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_434
timestamp 1607639953
transform 1 0 41014 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_422
timestamp 1607639953
transform 1 0 39910 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_459
timestamp 1607639953
transform 1 0 43314 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_446
timestamp 1607639953
transform 1 0 42118 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1607639953
transform 1 0 43222 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_483
timestamp 1607639953
transform 1 0 45522 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_471
timestamp 1607639953
transform 1 0 44418 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_495
timestamp 1607639953
transform 1 0 46626 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_520
timestamp 1607639953
transform 1 0 48926 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_507
timestamp 1607639953
transform 1 0 47730 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_722
timestamp 1607639953
transform 1 0 48834 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_544
timestamp 1607639953
transform 1 0 51134 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_532
timestamp 1607639953
transform 1 0 50030 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_568
timestamp 1607639953
transform 1 0 53342 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_556
timestamp 1607639953
transform 1 0 52238 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_593
timestamp 1607639953
transform 1 0 55642 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_581
timestamp 1607639953
transform 1 0 54538 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_723
timestamp 1607639953
transform 1 0 54446 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_605
timestamp 1607639953
transform 1 0 56746 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_617
timestamp 1607639953
transform 1 0 57850 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1607639953
transform -1 0 58862 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1607639953
transform 1 0 2466 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1607639953
transform 1 0 1362 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1607639953
transform 1 0 1086 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1607639953
transform 1 0 4674 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1607639953
transform 1 0 3570 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_62
timestamp 1607639953
transform 1 0 6790 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_59
timestamp 1607639953
transform 1 0 6514 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_51
timestamp 1607639953
transform 1 0 5778 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_724
timestamp 1607639953
transform 1 0 6698 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_74
timestamp 1607639953
transform 1 0 7894 0 1 29920
box -38 -48 222 592
use XNOR2X1  XNOR2X1
timestamp 1608122862
transform 1 0 8078 0 1 29920
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILLER_51_102
timestamp 1607639953
transform 1 0 10470 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_90
timestamp 1607639953
transform 1 0 9366 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_123
timestamp 1607639953
transform 1 0 12402 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_114
timestamp 1607639953
transform 1 0 11574 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_725
timestamp 1607639953
transform 1 0 12310 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_147
timestamp 1607639953
transform 1 0 14610 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_135
timestamp 1607639953
transform 1 0 13506 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_175
timestamp 1607639953
transform 1 0 17186 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_171
timestamp 1607639953
transform 1 0 16818 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_159
timestamp 1607639953
transform 1 0 15714 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1607639953
transform 1 0 16910 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_196
timestamp 1607639953
transform 1 0 19118 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_184
timestamp 1607639953
transform 1 0 18014 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_726
timestamp 1607639953
transform 1 0 17922 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_220
timestamp 1607639953
transform 1 0 21326 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_208
timestamp 1607639953
transform 1 0 20222 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_232
timestamp 1607639953
transform 1 0 22430 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_257
timestamp 1607639953
transform 1 0 24730 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_245
timestamp 1607639953
transform 1 0 23626 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_727
timestamp 1607639953
transform 1 0 23534 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1607639953
transform 1 0 26938 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_269
timestamp 1607639953
transform 1 0 25834 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1607639953
transform 1 0 28042 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_728
timestamp 1607639953
transform 1 0 29146 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _135_
timestamp 1607639953
transform 1 0 29238 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_321
timestamp 1607639953
transform 1 0 30618 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_309
timestamp 1607639953
transform 1 0 29514 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_345
timestamp 1607639953
transform 1 0 32826 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_333
timestamp 1607639953
transform 1 0 31722 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_367
timestamp 1607639953
transform 1 0 34850 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_365
timestamp 1607639953
transform 1 0 34666 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_357
timestamp 1607639953
transform 1 0 33930 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_729
timestamp 1607639953
transform 1 0 34758 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_391
timestamp 1607639953
transform 1 0 37058 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_379
timestamp 1607639953
transform 1 0 35954 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_415
timestamp 1607639953
transform 1 0 39266 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_403
timestamp 1607639953
transform 1 0 38162 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_440
timestamp 1607639953
transform 1 0 41566 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_428
timestamp 1607639953
transform 1 0 40462 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_730
timestamp 1607639953
transform 1 0 40370 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_452
timestamp 1607639953
transform 1 0 42670 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_476
timestamp 1607639953
transform 1 0 44878 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_464
timestamp 1607639953
transform 1 0 43774 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_501
timestamp 1607639953
transform 1 0 47178 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_489
timestamp 1607639953
transform 1 0 46074 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_731
timestamp 1607639953
transform 1 0 45982 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_528
timestamp 1607639953
transform 1 0 49662 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_516
timestamp 1607639953
transform 1 0 48558 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_512
timestamp 1607639953
transform 1 0 48190 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _173_
timestamp 1607639953
transform 1 0 48282 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1607639953
transform 1 0 47914 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_550
timestamp 1607639953
transform 1 0 51686 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_548
timestamp 1607639953
transform 1 0 51502 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_540
timestamp 1607639953
transform 1 0 50766 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_732
timestamp 1607639953
transform 1 0 51594 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_570
timestamp 1607639953
transform 1 0 53526 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_562
timestamp 1607639953
transform 1 0 52790 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_588
timestamp 1607639953
transform 1 0 55182 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_576
timestamp 1607639953
transform 1 0 54078 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _115_
timestamp 1607639953
transform 1 0 53802 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_611
timestamp 1607639953
transform 1 0 57298 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_608
timestamp 1607639953
transform 1 0 57022 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_600
timestamp 1607639953
transform 1 0 56286 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_733
timestamp 1607639953
transform 1 0 57206 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_623
timestamp 1607639953
transform 1 0 58402 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1607639953
transform -1 0 58862 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1607639953
transform 1 0 2466 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1607639953
transform 1 0 1362 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1607639953
transform 1 0 2466 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1607639953
transform 1 0 1362 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1607639953
transform 1 0 1086 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1607639953
transform 1 0 1086 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1607639953
transform 1 0 4674 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1607639953
transform 1 0 3570 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_44
timestamp 1607639953
transform 1 0 5134 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_32
timestamp 1607639953
transform 1 0 4030 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_27
timestamp 1607639953
transform 1 0 3570 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_734
timestamp 1607639953
transform 1 0 3938 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_62
timestamp 1607639953
transform 1 0 6790 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_59
timestamp 1607639953
transform 1 0 6514 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_51
timestamp 1607639953
transform 1 0 5778 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_56
timestamp 1607639953
transform 1 0 6238 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_744
timestamp 1607639953
transform 1 0 6698 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_74
timestamp 1607639953
transform 1 0 7894 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_80
timestamp 1607639953
transform 1 0 8446 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_68
timestamp 1607639953
transform 1 0 7342 0 -1 31008
box -38 -48 1142 592
use XOR2X1  XOR2X1
timestamp 1608122862
transform 1 0 8078 0 1 31008
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_6  FILLER_53_102
timestamp 1607639953
transform 1 0 10470 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_90
timestamp 1607639953
transform 1 0 9366 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_105
timestamp 1607639953
transform 1 0 10746 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_93
timestamp 1607639953
transform 1 0 9642 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_735
timestamp 1607639953
transform 1 0 9550 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _141_
timestamp 1607639953
transform 1 0 11022 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_123
timestamp 1607639953
transform 1 0 12402 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_119
timestamp 1607639953
transform 1 0 12034 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_111
timestamp 1607639953
transform 1 0 11298 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_129
timestamp 1607639953
transform 1 0 12954 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_117
timestamp 1607639953
transform 1 0 11850 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_745
timestamp 1607639953
transform 1 0 12310 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_147
timestamp 1607639953
transform 1 0 14610 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_135
timestamp 1607639953
transform 1 0 13506 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_154
timestamp 1607639953
transform 1 0 15254 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1607639953
transform 1 0 14058 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_736
timestamp 1607639953
transform 1 0 15162 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_171
timestamp 1607639953
transform 1 0 16818 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_159
timestamp 1607639953
transform 1 0 15714 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_166
timestamp 1607639953
transform 1 0 16358 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_196
timestamp 1607639953
transform 1 0 19118 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_184
timestamp 1607639953
transform 1 0 18014 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_190
timestamp 1607639953
transform 1 0 18566 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_178
timestamp 1607639953
transform 1 0 17462 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_746
timestamp 1607639953
transform 1 0 17922 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_220
timestamp 1607639953
transform 1 0 21326 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_208
timestamp 1607639953
transform 1 0 20222 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_215
timestamp 1607639953
transform 1 0 20866 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_202
timestamp 1607639953
transform 1 0 19670 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_737
timestamp 1607639953
transform 1 0 20774 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_232
timestamp 1607639953
transform 1 0 22430 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_239
timestamp 1607639953
transform 1 0 23074 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_227
timestamp 1607639953
transform 1 0 21970 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_257
timestamp 1607639953
transform 1 0 24730 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_245
timestamp 1607639953
transform 1 0 23626 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_263
timestamp 1607639953
transform 1 0 25282 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_251
timestamp 1607639953
transform 1 0 24178 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_747
timestamp 1607639953
transform 1 0 23534 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1607639953
transform 1 0 26938 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_269
timestamp 1607639953
transform 1 0 25834 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_276
timestamp 1607639953
transform 1 0 26478 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_738
timestamp 1607639953
transform 1 0 26386 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_306
timestamp 1607639953
transform 1 0 29238 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1607639953
transform 1 0 28042 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_300
timestamp 1607639953
transform 1 0 28686 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_288
timestamp 1607639953
transform 1 0 27582 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_748
timestamp 1607639953
transform 1 0 29146 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_330
timestamp 1607639953
transform 1 0 31446 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_318
timestamp 1607639953
transform 1 0 30342 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_324
timestamp 1607639953
transform 1 0 30894 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_312
timestamp 1607639953
transform 1 0 29790 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_342
timestamp 1607639953
transform 1 0 32550 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_349
timestamp 1607639953
transform 1 0 33194 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_337
timestamp 1607639953
transform 1 0 32090 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_739
timestamp 1607639953
transform 1 0 31998 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_367
timestamp 1607639953
transform 1 0 34850 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_354
timestamp 1607639953
transform 1 0 33654 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_373
timestamp 1607639953
transform 1 0 35402 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_361
timestamp 1607639953
transform 1 0 34298 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_749
timestamp 1607639953
transform 1 0 34758 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1607639953
transform 1 0 37242 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_381
timestamp 1607639953
transform 1 0 36138 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_375
timestamp 1607639953
transform 1 0 35586 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_385
timestamp 1607639953
transform 1 0 36506 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _118_
timestamp 1607639953
transform 1 0 35862 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_417
timestamp 1607639953
transform 1 0 39450 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1607639953
transform 1 0 38346 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_410
timestamp 1607639953
transform 1 0 38806 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_398
timestamp 1607639953
transform 1 0 37702 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_740
timestamp 1607639953
transform 1 0 37610 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_440
timestamp 1607639953
transform 1 0 41566 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_428
timestamp 1607639953
transform 1 0 40462 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_425
timestamp 1607639953
transform 1 0 40186 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_434
timestamp 1607639953
transform 1 0 41014 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_422
timestamp 1607639953
transform 1 0 39910 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_750
timestamp 1607639953
transform 1 0 40370 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_452
timestamp 1607639953
transform 1 0 42670 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_459
timestamp 1607639953
transform 1 0 43314 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_446
timestamp 1607639953
transform 1 0 42118 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_741
timestamp 1607639953
transform 1 0 43222 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_476
timestamp 1607639953
transform 1 0 44878 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_464
timestamp 1607639953
transform 1 0 43774 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_483
timestamp 1607639953
transform 1 0 45522 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_471
timestamp 1607639953
transform 1 0 44418 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_501
timestamp 1607639953
transform 1 0 47178 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_489
timestamp 1607639953
transform 1 0 46074 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_495
timestamp 1607639953
transform 1 0 46626 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_751
timestamp 1607639953
transform 1 0 45982 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_525
timestamp 1607639953
transform 1 0 49386 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_513
timestamp 1607639953
transform 1 0 48282 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_520
timestamp 1607639953
transform 1 0 48926 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_507
timestamp 1607639953
transform 1 0 47730 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_742
timestamp 1607639953
transform 1 0 48834 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_550
timestamp 1607639953
transform 1 0 51686 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_537
timestamp 1607639953
transform 1 0 50490 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_544
timestamp 1607639953
transform 1 0 51134 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_532
timestamp 1607639953
transform 1 0 50030 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_752
timestamp 1607639953
transform 1 0 51594 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_562
timestamp 1607639953
transform 1 0 52790 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_568
timestamp 1607639953
transform 1 0 53342 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_556
timestamp 1607639953
transform 1 0 52238 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_586
timestamp 1607639953
transform 1 0 54998 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_574
timestamp 1607639953
transform 1 0 53894 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_593
timestamp 1607639953
transform 1 0 55642 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_581
timestamp 1607639953
transform 1 0 54538 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_743
timestamp 1607639953
transform 1 0 54446 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_611
timestamp 1607639953
transform 1 0 57298 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_598
timestamp 1607639953
transform 1 0 56102 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_605
timestamp 1607639953
transform 1 0 56746 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_753
timestamp 1607639953
transform 1 0 57206 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_623
timestamp 1607639953
transform 1 0 58402 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_617
timestamp 1607639953
transform 1 0 57850 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1607639953
transform -1 0 58862 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1607639953
transform -1 0 58862 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1607639953
transform 1 0 2466 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1607639953
transform 1 0 1362 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1607639953
transform 1 0 1086 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_44
timestamp 1607639953
transform 1 0 5134 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_32
timestamp 1607639953
transform 1 0 4030 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_27
timestamp 1607639953
transform 1 0 3570 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_754
timestamp 1607639953
transform 1 0 3938 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_56
timestamp 1607639953
transform 1 0 6238 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_80
timestamp 1607639953
transform 1 0 8446 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_68
timestamp 1607639953
transform 1 0 7342 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_105
timestamp 1607639953
transform 1 0 10746 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_93
timestamp 1607639953
transform 1 0 9642 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_755
timestamp 1607639953
transform 1 0 9550 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_129
timestamp 1607639953
transform 1 0 12954 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_117
timestamp 1607639953
transform 1 0 11850 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_154
timestamp 1607639953
transform 1 0 15254 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1607639953
transform 1 0 14058 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_756
timestamp 1607639953
transform 1 0 15162 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_166
timestamp 1607639953
transform 1 0 16358 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_190
timestamp 1607639953
transform 1 0 18566 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_178
timestamp 1607639953
transform 1 0 17462 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_215
timestamp 1607639953
transform 1 0 20866 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_202
timestamp 1607639953
transform 1 0 19670 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_757
timestamp 1607639953
transform 1 0 20774 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_239
timestamp 1607639953
transform 1 0 23074 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_227
timestamp 1607639953
transform 1 0 21970 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_263
timestamp 1607639953
transform 1 0 25282 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_251
timestamp 1607639953
transform 1 0 24178 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_276
timestamp 1607639953
transform 1 0 26478 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_758
timestamp 1607639953
transform 1 0 26386 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_300
timestamp 1607639953
transform 1 0 28686 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_288
timestamp 1607639953
transform 1 0 27582 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_324
timestamp 1607639953
transform 1 0 30894 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_312
timestamp 1607639953
transform 1 0 29790 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_349
timestamp 1607639953
transform 1 0 33194 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_337
timestamp 1607639953
transform 1 0 32090 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_759
timestamp 1607639953
transform 1 0 31998 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_373
timestamp 1607639953
transform 1 0 35402 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_361
timestamp 1607639953
transform 1 0 34298 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_385
timestamp 1607639953
transform 1 0 36506 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_410
timestamp 1607639953
transform 1 0 38806 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_398
timestamp 1607639953
transform 1 0 37702 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_760
timestamp 1607639953
transform 1 0 37610 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_434
timestamp 1607639953
transform 1 0 41014 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_422
timestamp 1607639953
transform 1 0 39910 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_459
timestamp 1607639953
transform 1 0 43314 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_446
timestamp 1607639953
transform 1 0 42118 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_761
timestamp 1607639953
transform 1 0 43222 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_483
timestamp 1607639953
transform 1 0 45522 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_471
timestamp 1607639953
transform 1 0 44418 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_495
timestamp 1607639953
transform 1 0 46626 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_520
timestamp 1607639953
transform 1 0 48926 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_507
timestamp 1607639953
transform 1 0 47730 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_762
timestamp 1607639953
transform 1 0 48834 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_544
timestamp 1607639953
transform 1 0 51134 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_532
timestamp 1607639953
transform 1 0 50030 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_568
timestamp 1607639953
transform 1 0 53342 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_556
timestamp 1607639953
transform 1 0 52238 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_584
timestamp 1607639953
transform 1 0 54814 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_763
timestamp 1607639953
transform 1 0 54446 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _076_
timestamp 1607639953
transform 1 0 54538 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_608
timestamp 1607639953
transform 1 0 57022 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_596
timestamp 1607639953
transform 1 0 55918 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_624
timestamp 1607639953
transform 1 0 58494 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_620
timestamp 1607639953
transform 1 0 58126 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1607639953
transform -1 0 58862 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1607639953
transform 1 0 2466 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1607639953
transform 1 0 1362 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1607639953
transform 1 0 1086 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1607639953
transform 1 0 4674 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1607639953
transform 1 0 3570 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_62
timestamp 1607639953
transform 1 0 6790 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_59
timestamp 1607639953
transform 1 0 6514 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_51
timestamp 1607639953
transform 1 0 5778 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_764
timestamp 1607639953
transform 1 0 6698 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_86
timestamp 1607639953
transform 1 0 8998 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_74
timestamp 1607639953
transform 1 0 7894 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_110
timestamp 1607639953
transform 1 0 11206 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_98
timestamp 1607639953
transform 1 0 10102 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_123
timestamp 1607639953
transform 1 0 12402 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_765
timestamp 1607639953
transform 1 0 12310 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_147
timestamp 1607639953
transform 1 0 14610 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_135
timestamp 1607639953
transform 1 0 13506 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_171
timestamp 1607639953
transform 1 0 16818 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_159
timestamp 1607639953
transform 1 0 15714 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_196
timestamp 1607639953
transform 1 0 19118 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_184
timestamp 1607639953
transform 1 0 18014 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_766
timestamp 1607639953
transform 1 0 17922 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_220
timestamp 1607639953
transform 1 0 21326 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_208
timestamp 1607639953
transform 1 0 20222 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_232
timestamp 1607639953
transform 1 0 22430 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_257
timestamp 1607639953
transform 1 0 24730 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_245
timestamp 1607639953
transform 1 0 23626 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_767
timestamp 1607639953
transform 1 0 23534 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1607639953
transform 1 0 26938 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_269
timestamp 1607639953
transform 1 0 25834 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_306
timestamp 1607639953
transform 1 0 29238 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1607639953
transform 1 0 28042 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_768
timestamp 1607639953
transform 1 0 29146 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_330
timestamp 1607639953
transform 1 0 31446 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_318
timestamp 1607639953
transform 1 0 30342 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_342
timestamp 1607639953
transform 1 0 32550 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_367
timestamp 1607639953
transform 1 0 34850 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_354
timestamp 1607639953
transform 1 0 33654 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_769
timestamp 1607639953
transform 1 0 34758 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_391
timestamp 1607639953
transform 1 0 37058 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_379
timestamp 1607639953
transform 1 0 35954 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_415
timestamp 1607639953
transform 1 0 39266 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_403
timestamp 1607639953
transform 1 0 38162 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_440
timestamp 1607639953
transform 1 0 41566 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_428
timestamp 1607639953
transform 1 0 40462 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_770
timestamp 1607639953
transform 1 0 40370 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_452
timestamp 1607639953
transform 1 0 42670 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_476
timestamp 1607639953
transform 1 0 44878 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_464
timestamp 1607639953
transform 1 0 43774 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_501
timestamp 1607639953
transform 1 0 47178 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_489
timestamp 1607639953
transform 1 0 46074 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_771
timestamp 1607639953
transform 1 0 45982 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_525
timestamp 1607639953
transform 1 0 49386 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_513
timestamp 1607639953
transform 1 0 48282 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_550
timestamp 1607639953
transform 1 0 51686 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_537
timestamp 1607639953
transform 1 0 50490 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_772
timestamp 1607639953
transform 1 0 51594 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_562
timestamp 1607639953
transform 1 0 52790 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_586
timestamp 1607639953
transform 1 0 54998 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_574
timestamp 1607639953
transform 1 0 53894 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_611
timestamp 1607639953
transform 1 0 57298 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_598
timestamp 1607639953
transform 1 0 56102 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_773
timestamp 1607639953
transform 1 0 57206 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_623
timestamp 1607639953
transform 1 0 58402 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1607639953
transform -1 0 58862 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1607639953
transform 1 0 2466 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1607639953
transform 1 0 1362 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1607639953
transform 1 0 1086 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_36
timestamp 1607639953
transform 1 0 4398 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_32
timestamp 1607639953
transform 1 0 4030 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_27
timestamp 1607639953
transform 1 0 3570 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_774
timestamp 1607639953
transform 1 0 3938 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1607639953
transform 1 0 4122 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_60
timestamp 1607639953
transform 1 0 6606 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_48
timestamp 1607639953
transform 1 0 5502 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_84
timestamp 1607639953
transform 1 0 8814 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_72
timestamp 1607639953
transform 1 0 7710 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_105
timestamp 1607639953
transform 1 0 10746 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_93
timestamp 1607639953
transform 1 0 9642 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_775
timestamp 1607639953
transform 1 0 9550 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_130
timestamp 1607639953
transform 1 0 13046 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_118
timestamp 1607639953
transform 1 0 11942 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_113
timestamp 1607639953
transform 1 0 11482 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _177_
timestamp 1607639953
transform 1 0 11666 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_154
timestamp 1607639953
transform 1 0 15254 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_150
timestamp 1607639953
transform 1 0 14886 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_142
timestamp 1607639953
transform 1 0 14150 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_776
timestamp 1607639953
transform 1 0 15162 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_166
timestamp 1607639953
transform 1 0 16358 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_190
timestamp 1607639953
transform 1 0 18566 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_178
timestamp 1607639953
transform 1 0 17462 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_215
timestamp 1607639953
transform 1 0 20866 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_202
timestamp 1607639953
transform 1 0 19670 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_777
timestamp 1607639953
transform 1 0 20774 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_239
timestamp 1607639953
transform 1 0 23074 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_227
timestamp 1607639953
transform 1 0 21970 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_263
timestamp 1607639953
transform 1 0 25282 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_251
timestamp 1607639953
transform 1 0 24178 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_276
timestamp 1607639953
transform 1 0 26478 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_778
timestamp 1607639953
transform 1 0 26386 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_300
timestamp 1607639953
transform 1 0 28686 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_288
timestamp 1607639953
transform 1 0 27582 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_324
timestamp 1607639953
transform 1 0 30894 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_312
timestamp 1607639953
transform 1 0 29790 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_349
timestamp 1607639953
transform 1 0 33194 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_337
timestamp 1607639953
transform 1 0 32090 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_779
timestamp 1607639953
transform 1 0 31998 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_373
timestamp 1607639953
transform 1 0 35402 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_361
timestamp 1607639953
transform 1 0 34298 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_385
timestamp 1607639953
transform 1 0 36506 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_410
timestamp 1607639953
transform 1 0 38806 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_398
timestamp 1607639953
transform 1 0 37702 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_780
timestamp 1607639953
transform 1 0 37610 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_434
timestamp 1607639953
transform 1 0 41014 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_422
timestamp 1607639953
transform 1 0 39910 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_459
timestamp 1607639953
transform 1 0 43314 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_446
timestamp 1607639953
transform 1 0 42118 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_781
timestamp 1607639953
transform 1 0 43222 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_483
timestamp 1607639953
transform 1 0 45522 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_471
timestamp 1607639953
transform 1 0 44418 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_495
timestamp 1607639953
transform 1 0 46626 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_520
timestamp 1607639953
transform 1 0 48926 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_507
timestamp 1607639953
transform 1 0 47730 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_782
timestamp 1607639953
transform 1 0 48834 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_544
timestamp 1607639953
transform 1 0 51134 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_532
timestamp 1607639953
transform 1 0 50030 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_568
timestamp 1607639953
transform 1 0 53342 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_556
timestamp 1607639953
transform 1 0 52238 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_593
timestamp 1607639953
transform 1 0 55642 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_581
timestamp 1607639953
transform 1 0 54538 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_783
timestamp 1607639953
transform 1 0 54446 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_605
timestamp 1607639953
transform 1 0 56746 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_617
timestamp 1607639953
transform 1 0 57850 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1607639953
transform -1 0 58862 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1607639953
transform 1 0 2466 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1607639953
transform 1 0 1362 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1607639953
transform 1 0 1086 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1607639953
transform 1 0 4674 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1607639953
transform 1 0 3570 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_62
timestamp 1607639953
transform 1 0 6790 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_59
timestamp 1607639953
transform 1 0 6514 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_51
timestamp 1607639953
transform 1 0 5778 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_784
timestamp 1607639953
transform 1 0 6698 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_86
timestamp 1607639953
transform 1 0 8998 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_74
timestamp 1607639953
transform 1 0 7894 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_110
timestamp 1607639953
transform 1 0 11206 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_98
timestamp 1607639953
transform 1 0 10102 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_123
timestamp 1607639953
transform 1 0 12402 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_785
timestamp 1607639953
transform 1 0 12310 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_147
timestamp 1607639953
transform 1 0 14610 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_135
timestamp 1607639953
transform 1 0 13506 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_171
timestamp 1607639953
transform 1 0 16818 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_159
timestamp 1607639953
transform 1 0 15714 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_196
timestamp 1607639953
transform 1 0 19118 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_184
timestamp 1607639953
transform 1 0 18014 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_786
timestamp 1607639953
transform 1 0 17922 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_220
timestamp 1607639953
transform 1 0 21326 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_208
timestamp 1607639953
transform 1 0 20222 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_232
timestamp 1607639953
transform 1 0 22430 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_257
timestamp 1607639953
transform 1 0 24730 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_245
timestamp 1607639953
transform 1 0 23626 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_787
timestamp 1607639953
transform 1 0 23534 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1607639953
transform 1 0 26938 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_269
timestamp 1607639953
transform 1 0 25834 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_306
timestamp 1607639953
transform 1 0 29238 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1607639953
transform 1 0 28042 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_788
timestamp 1607639953
transform 1 0 29146 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_330
timestamp 1607639953
transform 1 0 31446 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_318
timestamp 1607639953
transform 1 0 30342 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_342
timestamp 1607639953
transform 1 0 32550 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_367
timestamp 1607639953
transform 1 0 34850 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_354
timestamp 1607639953
transform 1 0 33654 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_789
timestamp 1607639953
transform 1 0 34758 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_391
timestamp 1607639953
transform 1 0 37058 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_379
timestamp 1607639953
transform 1 0 35954 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_415
timestamp 1607639953
transform 1 0 39266 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_403
timestamp 1607639953
transform 1 0 38162 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_440
timestamp 1607639953
transform 1 0 41566 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_428
timestamp 1607639953
transform 1 0 40462 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_790
timestamp 1607639953
transform 1 0 40370 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_452
timestamp 1607639953
transform 1 0 42670 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_476
timestamp 1607639953
transform 1 0 44878 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_464
timestamp 1607639953
transform 1 0 43774 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_501
timestamp 1607639953
transform 1 0 47178 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_489
timestamp 1607639953
transform 1 0 46074 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_791
timestamp 1607639953
transform 1 0 45982 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_525
timestamp 1607639953
transform 1 0 49386 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_513
timestamp 1607639953
transform 1 0 48282 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_550
timestamp 1607639953
transform 1 0 51686 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_537
timestamp 1607639953
transform 1 0 50490 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_792
timestamp 1607639953
transform 1 0 51594 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_562
timestamp 1607639953
transform 1 0 52790 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_586
timestamp 1607639953
transform 1 0 54998 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_574
timestamp 1607639953
transform 1 0 53894 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_611
timestamp 1607639953
transform 1 0 57298 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_598
timestamp 1607639953
transform 1 0 56102 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_793
timestamp 1607639953
transform 1 0 57206 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_623
timestamp 1607639953
transform 1 0 58402 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1607639953
transform -1 0 58862 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1607639953
transform 1 0 2466 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1607639953
transform 1 0 1362 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1607639953
transform 1 0 1086 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_44
timestamp 1607639953
transform 1 0 5134 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_32
timestamp 1607639953
transform 1 0 4030 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_27
timestamp 1607639953
transform 1 0 3570 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_794
timestamp 1607639953
transform 1 0 3938 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_61
timestamp 1607639953
transform 1 0 6698 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_56
timestamp 1607639953
transform 1 0 6238 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _146_
timestamp 1607639953
transform 1 0 6422 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_85
timestamp 1607639953
transform 1 0 8906 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_73
timestamp 1607639953
transform 1 0 7802 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_105
timestamp 1607639953
transform 1 0 10746 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_93
timestamp 1607639953
transform 1 0 9642 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_91
timestamp 1607639953
transform 1 0 9458 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_795
timestamp 1607639953
transform 1 0 9550 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_129
timestamp 1607639953
transform 1 0 12954 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_117
timestamp 1607639953
transform 1 0 11850 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_154
timestamp 1607639953
transform 1 0 15254 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1607639953
transform 1 0 14058 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_796
timestamp 1607639953
transform 1 0 15162 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_166
timestamp 1607639953
transform 1 0 16358 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_190
timestamp 1607639953
transform 1 0 18566 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_178
timestamp 1607639953
transform 1 0 17462 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_215
timestamp 1607639953
transform 1 0 20866 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_202
timestamp 1607639953
transform 1 0 19670 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_797
timestamp 1607639953
transform 1 0 20774 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_239
timestamp 1607639953
transform 1 0 23074 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_227
timestamp 1607639953
transform 1 0 21970 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_263
timestamp 1607639953
transform 1 0 25282 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_251
timestamp 1607639953
transform 1 0 24178 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_276
timestamp 1607639953
transform 1 0 26478 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_798
timestamp 1607639953
transform 1 0 26386 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_300
timestamp 1607639953
transform 1 0 28686 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_288
timestamp 1607639953
transform 1 0 27582 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_324
timestamp 1607639953
transform 1 0 30894 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_312
timestamp 1607639953
transform 1 0 29790 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_349
timestamp 1607639953
transform 1 0 33194 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_337
timestamp 1607639953
transform 1 0 32090 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_799
timestamp 1607639953
transform 1 0 31998 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_373
timestamp 1607639953
transform 1 0 35402 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_361
timestamp 1607639953
transform 1 0 34298 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_385
timestamp 1607639953
transform 1 0 36506 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_410
timestamp 1607639953
transform 1 0 38806 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_398
timestamp 1607639953
transform 1 0 37702 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_800
timestamp 1607639953
transform 1 0 37610 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_434
timestamp 1607639953
transform 1 0 41014 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_422
timestamp 1607639953
transform 1 0 39910 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_459
timestamp 1607639953
transform 1 0 43314 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_446
timestamp 1607639953
transform 1 0 42118 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_801
timestamp 1607639953
transform 1 0 43222 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_483
timestamp 1607639953
transform 1 0 45522 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_471
timestamp 1607639953
transform 1 0 44418 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_495
timestamp 1607639953
transform 1 0 46626 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_520
timestamp 1607639953
transform 1 0 48926 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_507
timestamp 1607639953
transform 1 0 47730 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_802
timestamp 1607639953
transform 1 0 48834 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_544
timestamp 1607639953
transform 1 0 51134 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_532
timestamp 1607639953
transform 1 0 50030 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_568
timestamp 1607639953
transform 1 0 53342 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_556
timestamp 1607639953
transform 1 0 52238 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_593
timestamp 1607639953
transform 1 0 55642 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_581
timestamp 1607639953
transform 1 0 54538 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_803
timestamp 1607639953
transform 1 0 54446 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_605
timestamp 1607639953
transform 1 0 56746 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_617
timestamp 1607639953
transform 1 0 57850 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1607639953
transform -1 0 58862 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1607639953
transform 1 0 2466 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1607639953
transform 1 0 1362 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1607639953
transform 1 0 2466 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1607639953
transform 1 0 1362 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1607639953
transform 1 0 1086 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1607639953
transform 1 0 1086 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_44
timestamp 1607639953
transform 1 0 5134 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_32
timestamp 1607639953
transform 1 0 4030 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1607639953
transform 1 0 3570 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1607639953
transform 1 0 4674 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1607639953
transform 1 0 3570 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_814
timestamp 1607639953
transform 1 0 3938 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_56
timestamp 1607639953
transform 1 0 6238 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_62
timestamp 1607639953
transform 1 0 6790 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_59
timestamp 1607639953
transform 1 0 6514 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_51
timestamp 1607639953
transform 1 0 5778 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_804
timestamp 1607639953
transform 1 0 6698 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_80
timestamp 1607639953
transform 1 0 8446 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_68
timestamp 1607639953
transform 1 0 7342 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_86
timestamp 1607639953
transform 1 0 8998 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_74
timestamp 1607639953
transform 1 0 7894 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_105
timestamp 1607639953
transform 1 0 10746 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_93
timestamp 1607639953
transform 1 0 9642 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_110
timestamp 1607639953
transform 1 0 11206 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_98
timestamp 1607639953
transform 1 0 10102 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_815
timestamp 1607639953
transform 1 0 9550 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_129
timestamp 1607639953
transform 1 0 12954 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_117
timestamp 1607639953
transform 1 0 11850 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_123
timestamp 1607639953
transform 1 0 12402 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_805
timestamp 1607639953
transform 1 0 12310 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_154
timestamp 1607639953
transform 1 0 15254 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1607639953
transform 1 0 14058 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_147
timestamp 1607639953
transform 1 0 14610 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_135
timestamp 1607639953
transform 1 0 13506 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_816
timestamp 1607639953
transform 1 0 15162 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_166
timestamp 1607639953
transform 1 0 16358 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_162
timestamp 1607639953
transform 1 0 15990 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_171
timestamp 1607639953
transform 1 0 16818 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_159
timestamp 1607639953
transform 1 0 15714 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _174_
timestamp 1607639953
transform 1 0 16082 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_190
timestamp 1607639953
transform 1 0 18566 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_178
timestamp 1607639953
transform 1 0 17462 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_196
timestamp 1607639953
transform 1 0 19118 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_184
timestamp 1607639953
transform 1 0 18014 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_806
timestamp 1607639953
transform 1 0 17922 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_215
timestamp 1607639953
transform 1 0 20866 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_202
timestamp 1607639953
transform 1 0 19670 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_220
timestamp 1607639953
transform 1 0 21326 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_208
timestamp 1607639953
transform 1 0 20222 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_817
timestamp 1607639953
transform 1 0 20774 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_239
timestamp 1607639953
transform 1 0 23074 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_227
timestamp 1607639953
transform 1 0 21970 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_232
timestamp 1607639953
transform 1 0 22430 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_263
timestamp 1607639953
transform 1 0 25282 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_251
timestamp 1607639953
transform 1 0 24178 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_257
timestamp 1607639953
transform 1 0 24730 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_245
timestamp 1607639953
transform 1 0 23626 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_807
timestamp 1607639953
transform 1 0 23534 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_276
timestamp 1607639953
transform 1 0 26478 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1607639953
transform 1 0 26938 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_269
timestamp 1607639953
transform 1 0 25834 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_818
timestamp 1607639953
transform 1 0 26386 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_300
timestamp 1607639953
transform 1 0 28686 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_288
timestamp 1607639953
transform 1 0 27582 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_306
timestamp 1607639953
transform 1 0 29238 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1607639953
transform 1 0 28042 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_808
timestamp 1607639953
transform 1 0 29146 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_324
timestamp 1607639953
transform 1 0 30894 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_312
timestamp 1607639953
transform 1 0 29790 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_330
timestamp 1607639953
transform 1 0 31446 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_318
timestamp 1607639953
transform 1 0 30342 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_349
timestamp 1607639953
transform 1 0 33194 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_337
timestamp 1607639953
transform 1 0 32090 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_342
timestamp 1607639953
transform 1 0 32550 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_819
timestamp 1607639953
transform 1 0 31998 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_373
timestamp 1607639953
transform 1 0 35402 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_361
timestamp 1607639953
transform 1 0 34298 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_367
timestamp 1607639953
transform 1 0 34850 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_354
timestamp 1607639953
transform 1 0 33654 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_809
timestamp 1607639953
transform 1 0 34758 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_385
timestamp 1607639953
transform 1 0 36506 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_391
timestamp 1607639953
transform 1 0 37058 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_379
timestamp 1607639953
transform 1 0 35954 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_410
timestamp 1607639953
transform 1 0 38806 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_398
timestamp 1607639953
transform 1 0 37702 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_415
timestamp 1607639953
transform 1 0 39266 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_403
timestamp 1607639953
transform 1 0 38162 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_820
timestamp 1607639953
transform 1 0 37610 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_434
timestamp 1607639953
transform 1 0 41014 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_422
timestamp 1607639953
transform 1 0 39910 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_440
timestamp 1607639953
transform 1 0 41566 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_428
timestamp 1607639953
transform 1 0 40462 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_810
timestamp 1607639953
transform 1 0 40370 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_459
timestamp 1607639953
transform 1 0 43314 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_446
timestamp 1607639953
transform 1 0 42118 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_457
timestamp 1607639953
transform 1 0 43130 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_452
timestamp 1607639953
transform 1 0 42670 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_821
timestamp 1607639953
transform 1 0 43222 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _132_
timestamp 1607639953
transform 1 0 42854 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_483
timestamp 1607639953
transform 1 0 45522 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_471
timestamp 1607639953
transform 1 0 44418 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_481
timestamp 1607639953
transform 1 0 45338 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_469
timestamp 1607639953
transform 1 0 44234 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_495
timestamp 1607639953
transform 1 0 46626 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_501
timestamp 1607639953
transform 1 0 47178 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_489
timestamp 1607639953
transform 1 0 46074 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_487
timestamp 1607639953
transform 1 0 45890 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_811
timestamp 1607639953
transform 1 0 45982 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_520
timestamp 1607639953
transform 1 0 48926 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_507
timestamp 1607639953
transform 1 0 47730 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_525
timestamp 1607639953
transform 1 0 49386 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_513
timestamp 1607639953
transform 1 0 48282 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_822
timestamp 1607639953
transform 1 0 48834 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_544
timestamp 1607639953
transform 1 0 51134 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_532
timestamp 1607639953
transform 1 0 50030 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_550
timestamp 1607639953
transform 1 0 51686 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_537
timestamp 1607639953
transform 1 0 50490 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_812
timestamp 1607639953
transform 1 0 51594 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_568
timestamp 1607639953
transform 1 0 53342 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_556
timestamp 1607639953
transform 1 0 52238 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_562
timestamp 1607639953
transform 1 0 52790 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_593
timestamp 1607639953
transform 1 0 55642 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_581
timestamp 1607639953
transform 1 0 54538 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_586
timestamp 1607639953
transform 1 0 54998 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_574
timestamp 1607639953
transform 1 0 53894 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_823
timestamp 1607639953
transform 1 0 54446 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_605
timestamp 1607639953
transform 1 0 56746 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_611
timestamp 1607639953
transform 1 0 57298 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_598
timestamp 1607639953
transform 1 0 56102 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_813
timestamp 1607639953
transform 1 0 57206 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_617
timestamp 1607639953
transform 1 0 57850 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_623
timestamp 1607639953
transform 1 0 58402 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1607639953
transform -1 0 58862 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1607639953
transform -1 0 58862 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1607639953
transform 1 0 2466 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1607639953
transform 1 0 1362 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1607639953
transform 1 0 1086 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_38
timestamp 1607639953
transform 1 0 4582 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_27
timestamp 1607639953
transform 1 0 3570 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _079_
timestamp 1607639953
transform 1 0 4306 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_62
timestamp 1607639953
transform 1 0 6790 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_58
timestamp 1607639953
transform 1 0 6422 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_50
timestamp 1607639953
transform 1 0 5686 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_824
timestamp 1607639953
transform 1 0 6698 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_86
timestamp 1607639953
transform 1 0 8998 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_74
timestamp 1607639953
transform 1 0 7894 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_110
timestamp 1607639953
transform 1 0 11206 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_98
timestamp 1607639953
transform 1 0 10102 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_123
timestamp 1607639953
transform 1 0 12402 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_825
timestamp 1607639953
transform 1 0 12310 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_147
timestamp 1607639953
transform 1 0 14610 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_135
timestamp 1607639953
transform 1 0 13506 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_171
timestamp 1607639953
transform 1 0 16818 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_159
timestamp 1607639953
transform 1 0 15714 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_196
timestamp 1607639953
transform 1 0 19118 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_184
timestamp 1607639953
transform 1 0 18014 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_826
timestamp 1607639953
transform 1 0 17922 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_220
timestamp 1607639953
transform 1 0 21326 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_208
timestamp 1607639953
transform 1 0 20222 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_232
timestamp 1607639953
transform 1 0 22430 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_257
timestamp 1607639953
transform 1 0 24730 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_245
timestamp 1607639953
transform 1 0 23626 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_827
timestamp 1607639953
transform 1 0 23534 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1607639953
transform 1 0 26938 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_269
timestamp 1607639953
transform 1 0 25834 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_306
timestamp 1607639953
transform 1 0 29238 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1607639953
transform 1 0 28042 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_828
timestamp 1607639953
transform 1 0 29146 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_330
timestamp 1607639953
transform 1 0 31446 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_318
timestamp 1607639953
transform 1 0 30342 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_342
timestamp 1607639953
transform 1 0 32550 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_367
timestamp 1607639953
transform 1 0 34850 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_354
timestamp 1607639953
transform 1 0 33654 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_829
timestamp 1607639953
transform 1 0 34758 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_391
timestamp 1607639953
transform 1 0 37058 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_379
timestamp 1607639953
transform 1 0 35954 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_418
timestamp 1607639953
transform 1 0 39542 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_406
timestamp 1607639953
transform 1 0 38438 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1607639953
transform 1 0 38162 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_440
timestamp 1607639953
transform 1 0 41566 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_428
timestamp 1607639953
transform 1 0 40462 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_426
timestamp 1607639953
transform 1 0 40278 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_830
timestamp 1607639953
transform 1 0 40370 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_452
timestamp 1607639953
transform 1 0 42670 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_476
timestamp 1607639953
transform 1 0 44878 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_464
timestamp 1607639953
transform 1 0 43774 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_501
timestamp 1607639953
transform 1 0 47178 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_489
timestamp 1607639953
transform 1 0 46074 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_831
timestamp 1607639953
transform 1 0 45982 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_525
timestamp 1607639953
transform 1 0 49386 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_513
timestamp 1607639953
transform 1 0 48282 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_550
timestamp 1607639953
transform 1 0 51686 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_537
timestamp 1607639953
transform 1 0 50490 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_832
timestamp 1607639953
transform 1 0 51594 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_562
timestamp 1607639953
transform 1 0 52790 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_594
timestamp 1607639953
transform 1 0 55734 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_590
timestamp 1607639953
transform 1 0 55366 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_586
timestamp 1607639953
transform 1 0 54998 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_574
timestamp 1607639953
transform 1 0 53894 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _162_
timestamp 1607639953
transform 1 0 55458 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_611
timestamp 1607639953
transform 1 0 57298 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_606
timestamp 1607639953
transform 1 0 56838 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_833
timestamp 1607639953
transform 1 0 57206 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_623
timestamp 1607639953
transform 1 0 58402 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1607639953
transform -1 0 58862 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1607639953
transform 1 0 2466 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1607639953
transform 1 0 1362 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1607639953
transform 1 0 1086 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_44
timestamp 1607639953
transform 1 0 5134 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_32
timestamp 1607639953
transform 1 0 4030 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1607639953
transform 1 0 3570 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_834
timestamp 1607639953
transform 1 0 3938 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_58
timestamp 1607639953
transform 1 0 6422 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_52
timestamp 1607639953
transform 1 0 5870 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _107_
timestamp 1607639953
transform 1 0 6146 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_82
timestamp 1607639953
transform 1 0 8630 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_70
timestamp 1607639953
transform 1 0 7526 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_105
timestamp 1607639953
transform 1 0 10746 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_93
timestamp 1607639953
transform 1 0 9642 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_90
timestamp 1607639953
transform 1 0 9366 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_835
timestamp 1607639953
transform 1 0 9550 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_129
timestamp 1607639953
transform 1 0 12954 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_117
timestamp 1607639953
transform 1 0 11850 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_154
timestamp 1607639953
transform 1 0 15254 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1607639953
transform 1 0 14058 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_836
timestamp 1607639953
transform 1 0 15162 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_166
timestamp 1607639953
transform 1 0 16358 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_190
timestamp 1607639953
transform 1 0 18566 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_178
timestamp 1607639953
transform 1 0 17462 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_215
timestamp 1607639953
transform 1 0 20866 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_202
timestamp 1607639953
transform 1 0 19670 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_837
timestamp 1607639953
transform 1 0 20774 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_239
timestamp 1607639953
transform 1 0 23074 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_227
timestamp 1607639953
transform 1 0 21970 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_263
timestamp 1607639953
transform 1 0 25282 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_251
timestamp 1607639953
transform 1 0 24178 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_276
timestamp 1607639953
transform 1 0 26478 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_838
timestamp 1607639953
transform 1 0 26386 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_300
timestamp 1607639953
transform 1 0 28686 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_288
timestamp 1607639953
transform 1 0 27582 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_324
timestamp 1607639953
transform 1 0 30894 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_312
timestamp 1607639953
transform 1 0 29790 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_349
timestamp 1607639953
transform 1 0 33194 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_337
timestamp 1607639953
transform 1 0 32090 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_839
timestamp 1607639953
transform 1 0 31998 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_373
timestamp 1607639953
transform 1 0 35402 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_361
timestamp 1607639953
transform 1 0 34298 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_385
timestamp 1607639953
transform 1 0 36506 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_415
timestamp 1607639953
transform 1 0 39266 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_403
timestamp 1607639953
transform 1 0 38162 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_398
timestamp 1607639953
transform 1 0 37702 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_840
timestamp 1607639953
transform 1 0 37610 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _140_
timestamp 1607639953
transform 1 0 37886 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_439
timestamp 1607639953
transform 1 0 41474 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_427
timestamp 1607639953
transform 1 0 40370 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_459
timestamp 1607639953
transform 1 0 43314 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_457
timestamp 1607639953
transform 1 0 43130 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_451
timestamp 1607639953
transform 1 0 42578 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_841
timestamp 1607639953
transform 1 0 43222 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_483
timestamp 1607639953
transform 1 0 45522 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_471
timestamp 1607639953
transform 1 0 44418 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_495
timestamp 1607639953
transform 1 0 46626 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_520
timestamp 1607639953
transform 1 0 48926 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_507
timestamp 1607639953
transform 1 0 47730 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_842
timestamp 1607639953
transform 1 0 48834 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_544
timestamp 1607639953
transform 1 0 51134 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_532
timestamp 1607639953
transform 1 0 50030 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_568
timestamp 1607639953
transform 1 0 53342 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_556
timestamp 1607639953
transform 1 0 52238 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_593
timestamp 1607639953
transform 1 0 55642 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_581
timestamp 1607639953
transform 1 0 54538 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_843
timestamp 1607639953
transform 1 0 54446 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_605
timestamp 1607639953
transform 1 0 56746 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_617
timestamp 1607639953
transform 1 0 57850 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1607639953
transform -1 0 58862 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1607639953
transform 1 0 2466 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1607639953
transform 1 0 1362 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1607639953
transform 1 0 1086 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_40
timestamp 1607639953
transform 1 0 4766 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_35
timestamp 1607639953
transform 1 0 4306 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_27
timestamp 1607639953
transform 1 0 3570 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _180_
timestamp 1607639953
transform 1 0 4490 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_62
timestamp 1607639953
transform 1 0 6790 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_60
timestamp 1607639953
transform 1 0 6606 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_52
timestamp 1607639953
transform 1 0 5870 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_844
timestamp 1607639953
transform 1 0 6698 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_86
timestamp 1607639953
transform 1 0 8998 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_74
timestamp 1607639953
transform 1 0 7894 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_110
timestamp 1607639953
transform 1 0 11206 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_98
timestamp 1607639953
transform 1 0 10102 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1607639953
transform 1 0 12402 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_121
timestamp 1607639953
transform 1 0 12218 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_117
timestamp 1607639953
transform 1 0 11850 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_845
timestamp 1607639953
transform 1 0 12310 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _193_
timestamp 1607639953
transform 1 0 11574 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_63_153
timestamp 1607639953
transform 1 0 15162 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_147
timestamp 1607639953
transform 1 0 14610 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_135
timestamp 1607639953
transform 1 0 13506 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _150_
timestamp 1607639953
transform 1 0 15254 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1607639953
transform 1 0 16634 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_157
timestamp 1607639953
transform 1 0 15530 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_196
timestamp 1607639953
transform 1 0 19118 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_184
timestamp 1607639953
transform 1 0 18014 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_181
timestamp 1607639953
transform 1 0 17738 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_846
timestamp 1607639953
transform 1 0 17922 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1607639953
transform 1 0 19210 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_212
timestamp 1607639953
transform 1 0 20590 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_200
timestamp 1607639953
transform 1 0 19486 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_236
timestamp 1607639953
transform 1 0 22798 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_224
timestamp 1607639953
transform 1 0 21694 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_257
timestamp 1607639953
transform 1 0 24730 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_245
timestamp 1607639953
transform 1 0 23626 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_847
timestamp 1607639953
transform 1 0 23534 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1607639953
transform 1 0 26938 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_269
timestamp 1607639953
transform 1 0 25834 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_306
timestamp 1607639953
transform 1 0 29238 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1607639953
transform 1 0 28042 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_848
timestamp 1607639953
transform 1 0 29146 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_330
timestamp 1607639953
transform 1 0 31446 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_318
timestamp 1607639953
transform 1 0 30342 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_342
timestamp 1607639953
transform 1 0 32550 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_370
timestamp 1607639953
transform 1 0 35126 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_354
timestamp 1607639953
transform 1 0 33654 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_849
timestamp 1607639953
transform 1 0 34758 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _123_
timestamp 1607639953
transform 1 0 34850 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_394
timestamp 1607639953
transform 1 0 37334 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_382
timestamp 1607639953
transform 1 0 36230 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_418
timestamp 1607639953
transform 1 0 39542 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_406
timestamp 1607639953
transform 1 0 38438 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_440
timestamp 1607639953
transform 1 0 41566 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_428
timestamp 1607639953
transform 1 0 40462 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_426
timestamp 1607639953
transform 1 0 40278 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_850
timestamp 1607639953
transform 1 0 40370 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_452
timestamp 1607639953
transform 1 0 42670 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_476
timestamp 1607639953
transform 1 0 44878 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_464
timestamp 1607639953
transform 1 0 43774 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_501
timestamp 1607639953
transform 1 0 47178 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_489
timestamp 1607639953
transform 1 0 46074 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_851
timestamp 1607639953
transform 1 0 45982 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_525
timestamp 1607639953
transform 1 0 49386 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_513
timestamp 1607639953
transform 1 0 48282 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_550
timestamp 1607639953
transform 1 0 51686 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_537
timestamp 1607639953
transform 1 0 50490 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_852
timestamp 1607639953
transform 1 0 51594 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_566
timestamp 1607639953
transform 1 0 53158 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_562
timestamp 1607639953
transform 1 0 52790 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1607639953
transform 1 0 52882 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_590
timestamp 1607639953
transform 1 0 55366 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_578
timestamp 1607639953
transform 1 0 54262 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_611
timestamp 1607639953
transform 1 0 57298 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_602
timestamp 1607639953
transform 1 0 56470 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_853
timestamp 1607639953
transform 1 0 57206 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_623
timestamp 1607639953
transform 1 0 58402 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1607639953
transform -1 0 58862 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1607639953
transform 1 0 2466 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1607639953
transform 1 0 1362 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1607639953
transform 1 0 1086 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_44
timestamp 1607639953
transform 1 0 5134 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1607639953
transform 1 0 4030 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1607639953
transform 1 0 3570 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_854
timestamp 1607639953
transform 1 0 3938 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_56
timestamp 1607639953
transform 1 0 6238 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_80
timestamp 1607639953
transform 1 0 8446 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_68
timestamp 1607639953
transform 1 0 7342 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_110
timestamp 1607639953
transform 1 0 11206 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_105
timestamp 1607639953
transform 1 0 10746 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_93
timestamp 1607639953
transform 1 0 9642 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_855
timestamp 1607639953
transform 1 0 9550 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _138_
timestamp 1607639953
transform 1 0 10930 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_122
timestamp 1607639953
transform 1 0 12310 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_154
timestamp 1607639953
transform 1 0 15254 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_152
timestamp 1607639953
transform 1 0 15070 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_146
timestamp 1607639953
transform 1 0 14518 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_134
timestamp 1607639953
transform 1 0 13414 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_856
timestamp 1607639953
transform 1 0 15162 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_166
timestamp 1607639953
transform 1 0 16358 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_190
timestamp 1607639953
transform 1 0 18566 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_178
timestamp 1607639953
transform 1 0 17462 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_215
timestamp 1607639953
transform 1 0 20866 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_202
timestamp 1607639953
transform 1 0 19670 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_857
timestamp 1607639953
transform 1 0 20774 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_240
timestamp 1607639953
transform 1 0 23166 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_228
timestamp 1607639953
transform 1 0 22062 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_223
timestamp 1607639953
transform 1 0 21602 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _005_
timestamp 1607639953
transform 1 0 21786 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_264
timestamp 1607639953
transform 1 0 25374 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_260
timestamp 1607639953
transform 1 0 25006 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_252
timestamp 1607639953
transform 1 0 24270 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1607639953
transform 1 0 25098 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_282
timestamp 1607639953
transform 1 0 27030 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_276
timestamp 1607639953
transform 1 0 26478 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_272
timestamp 1607639953
transform 1 0 26110 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_858
timestamp 1607639953
transform 1 0 26386 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1607639953
transform 1 0 26754 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_306
timestamp 1607639953
transform 1 0 29238 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_294
timestamp 1607639953
transform 1 0 28134 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_330
timestamp 1607639953
transform 1 0 31446 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_318
timestamp 1607639953
transform 1 0 30342 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_349
timestamp 1607639953
transform 1 0 33194 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_337
timestamp 1607639953
transform 1 0 32090 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_859
timestamp 1607639953
transform 1 0 31998 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_373
timestamp 1607639953
transform 1 0 35402 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_361
timestamp 1607639953
transform 1 0 34298 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_385
timestamp 1607639953
transform 1 0 36506 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_410
timestamp 1607639953
transform 1 0 38806 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_398
timestamp 1607639953
transform 1 0 37702 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_860
timestamp 1607639953
transform 1 0 37610 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_434
timestamp 1607639953
transform 1 0 41014 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_422
timestamp 1607639953
transform 1 0 39910 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_459
timestamp 1607639953
transform 1 0 43314 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_446
timestamp 1607639953
transform 1 0 42118 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_861
timestamp 1607639953
transform 1 0 43222 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_479
timestamp 1607639953
transform 1 0 45154 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1607639953
transform 1 0 44786 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_471
timestamp 1607639953
transform 1 0 44418 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _113_
timestamp 1607639953
transform 1 0 44878 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_503
timestamp 1607639953
transform 1 0 47362 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_491
timestamp 1607639953
transform 1 0 46258 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_520
timestamp 1607639953
transform 1 0 48926 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_515
timestamp 1607639953
transform 1 0 48466 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_862
timestamp 1607639953
transform 1 0 48834 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_544
timestamp 1607639953
transform 1 0 51134 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_532
timestamp 1607639953
transform 1 0 50030 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_568
timestamp 1607639953
transform 1 0 53342 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_556
timestamp 1607639953
transform 1 0 52238 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_593
timestamp 1607639953
transform 1 0 55642 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_581
timestamp 1607639953
transform 1 0 54538 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_863
timestamp 1607639953
transform 1 0 54446 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_605
timestamp 1607639953
transform 1 0 56746 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_617
timestamp 1607639953
transform 1 0 57850 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1607639953
transform -1 0 58862 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1607639953
transform 1 0 2466 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1607639953
transform 1 0 1362 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1607639953
transform 1 0 1086 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1607639953
transform 1 0 4674 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1607639953
transform 1 0 3570 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_62
timestamp 1607639953
transform 1 0 6790 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_59
timestamp 1607639953
transform 1 0 6514 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_51
timestamp 1607639953
transform 1 0 5778 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_864
timestamp 1607639953
transform 1 0 6698 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_86
timestamp 1607639953
transform 1 0 8998 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_74
timestamp 1607639953
transform 1 0 7894 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_110
timestamp 1607639953
transform 1 0 11206 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_98
timestamp 1607639953
transform 1 0 10102 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_123
timestamp 1607639953
transform 1 0 12402 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_865
timestamp 1607639953
transform 1 0 12310 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_147
timestamp 1607639953
transform 1 0 14610 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_135
timestamp 1607639953
transform 1 0 13506 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_171
timestamp 1607639953
transform 1 0 16818 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_159
timestamp 1607639953
transform 1 0 15714 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_196
timestamp 1607639953
transform 1 0 19118 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_184
timestamp 1607639953
transform 1 0 18014 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_866
timestamp 1607639953
transform 1 0 17922 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_220
timestamp 1607639953
transform 1 0 21326 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_208
timestamp 1607639953
transform 1 0 20222 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_232
timestamp 1607639953
transform 1 0 22430 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_257
timestamp 1607639953
transform 1 0 24730 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_245
timestamp 1607639953
transform 1 0 23626 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_867
timestamp 1607639953
transform 1 0 23534 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1607639953
transform 1 0 26938 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_269
timestamp 1607639953
transform 1 0 25834 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_306
timestamp 1607639953
transform 1 0 29238 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1607639953
transform 1 0 28042 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_868
timestamp 1607639953
transform 1 0 29146 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_330
timestamp 1607639953
transform 1 0 31446 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_318
timestamp 1607639953
transform 1 0 30342 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_342
timestamp 1607639953
transform 1 0 32550 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_367
timestamp 1607639953
transform 1 0 34850 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_354
timestamp 1607639953
transform 1 0 33654 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_869
timestamp 1607639953
transform 1 0 34758 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_391
timestamp 1607639953
transform 1 0 37058 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_379
timestamp 1607639953
transform 1 0 35954 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_415
timestamp 1607639953
transform 1 0 39266 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_403
timestamp 1607639953
transform 1 0 38162 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_440
timestamp 1607639953
transform 1 0 41566 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_428
timestamp 1607639953
transform 1 0 40462 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_870
timestamp 1607639953
transform 1 0 40370 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_452
timestamp 1607639953
transform 1 0 42670 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_476
timestamp 1607639953
transform 1 0 44878 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_464
timestamp 1607639953
transform 1 0 43774 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_501
timestamp 1607639953
transform 1 0 47178 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_489
timestamp 1607639953
transform 1 0 46074 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_871
timestamp 1607639953
transform 1 0 45982 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_525
timestamp 1607639953
transform 1 0 49386 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_513
timestamp 1607639953
transform 1 0 48282 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_550
timestamp 1607639953
transform 1 0 51686 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_537
timestamp 1607639953
transform 1 0 50490 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_872
timestamp 1607639953
transform 1 0 51594 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_562
timestamp 1607639953
transform 1 0 52790 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_586
timestamp 1607639953
transform 1 0 54998 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_574
timestamp 1607639953
transform 1 0 53894 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_611
timestamp 1607639953
transform 1 0 57298 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_598
timestamp 1607639953
transform 1 0 56102 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_873
timestamp 1607639953
transform 1 0 57206 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_623
timestamp 1607639953
transform 1 0 58402 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1607639953
transform -1 0 58862 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1607639953
transform 1 0 2466 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1607639953
transform 1 0 1362 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1607639953
transform 1 0 2466 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1607639953
transform 1 0 1362 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1607639953
transform 1 0 1086 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1607639953
transform 1 0 1086 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1607639953
transform 1 0 4674 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1607639953
transform 1 0 3570 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_44
timestamp 1607639953
transform 1 0 5134 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_32
timestamp 1607639953
transform 1 0 4030 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_27
timestamp 1607639953
transform 1 0 3570 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_874
timestamp 1607639953
transform 1 0 3938 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_62
timestamp 1607639953
transform 1 0 6790 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_59
timestamp 1607639953
transform 1 0 6514 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_51
timestamp 1607639953
transform 1 0 5778 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_56
timestamp 1607639953
transform 1 0 6238 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_884
timestamp 1607639953
transform 1 0 6698 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_86
timestamp 1607639953
transform 1 0 8998 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_74
timestamp 1607639953
transform 1 0 7894 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_80
timestamp 1607639953
transform 1 0 8446 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_68
timestamp 1607639953
transform 1 0 7342 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_110
timestamp 1607639953
transform 1 0 11206 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_98
timestamp 1607639953
transform 1 0 10102 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_105
timestamp 1607639953
transform 1 0 10746 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_93
timestamp 1607639953
transform 1 0 9642 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_875
timestamp 1607639953
transform 1 0 9550 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_123
timestamp 1607639953
transform 1 0 12402 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_129
timestamp 1607639953
transform 1 0 12954 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_117
timestamp 1607639953
transform 1 0 11850 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_885
timestamp 1607639953
transform 1 0 12310 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_147
timestamp 1607639953
transform 1 0 14610 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_135
timestamp 1607639953
transform 1 0 13506 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_154
timestamp 1607639953
transform 1 0 15254 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1607639953
transform 1 0 14058 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_876
timestamp 1607639953
transform 1 0 15162 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_171
timestamp 1607639953
transform 1 0 16818 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_159
timestamp 1607639953
transform 1 0 15714 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_166
timestamp 1607639953
transform 1 0 16358 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_196
timestamp 1607639953
transform 1 0 19118 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_184
timestamp 1607639953
transform 1 0 18014 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_190
timestamp 1607639953
transform 1 0 18566 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_178
timestamp 1607639953
transform 1 0 17462 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_886
timestamp 1607639953
transform 1 0 17922 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_220
timestamp 1607639953
transform 1 0 21326 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_208
timestamp 1607639953
transform 1 0 20222 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_215
timestamp 1607639953
transform 1 0 20866 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_202
timestamp 1607639953
transform 1 0 19670 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_877
timestamp 1607639953
transform 1 0 20774 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_241
timestamp 1607639953
transform 1 0 23258 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_232
timestamp 1607639953
transform 1 0 22430 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_239
timestamp 1607639953
transform 1 0 23074 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_227
timestamp 1607639953
transform 1 0 21970 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1607639953
transform 1 0 22982 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_257
timestamp 1607639953
transform 1 0 24730 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_245
timestamp 1607639953
transform 1 0 23626 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_263
timestamp 1607639953
transform 1 0 25282 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_251
timestamp 1607639953
transform 1 0 24178 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_887
timestamp 1607639953
transform 1 0 23534 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1607639953
transform 1 0 26938 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_269
timestamp 1607639953
transform 1 0 25834 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_279
timestamp 1607639953
transform 1 0 26754 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_878
timestamp 1607639953
transform 1 0 26386 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _091_
timestamp 1607639953
transform 1 0 26478 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_306
timestamp 1607639953
transform 1 0 29238 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1607639953
transform 1 0 28042 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_303
timestamp 1607639953
transform 1 0 28962 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_291
timestamp 1607639953
transform 1 0 27858 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_888
timestamp 1607639953
transform 1 0 29146 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_330
timestamp 1607639953
transform 1 0 31446 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_318
timestamp 1607639953
transform 1 0 30342 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_327
timestamp 1607639953
transform 1 0 31170 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_315
timestamp 1607639953
transform 1 0 30066 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_342
timestamp 1607639953
transform 1 0 32550 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_349
timestamp 1607639953
transform 1 0 33194 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_337
timestamp 1607639953
transform 1 0 32090 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_335
timestamp 1607639953
transform 1 0 31906 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_879
timestamp 1607639953
transform 1 0 31998 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_367
timestamp 1607639953
transform 1 0 34850 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_354
timestamp 1607639953
transform 1 0 33654 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_373
timestamp 1607639953
transform 1 0 35402 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_361
timestamp 1607639953
transform 1 0 34298 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_889
timestamp 1607639953
transform 1 0 34758 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_391
timestamp 1607639953
transform 1 0 37058 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_379
timestamp 1607639953
transform 1 0 35954 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_385
timestamp 1607639953
transform 1 0 36506 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_415
timestamp 1607639953
transform 1 0 39266 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_403
timestamp 1607639953
transform 1 0 38162 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_410
timestamp 1607639953
transform 1 0 38806 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_398
timestamp 1607639953
transform 1 0 37702 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_880
timestamp 1607639953
transform 1 0 37610 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_440
timestamp 1607639953
transform 1 0 41566 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_428
timestamp 1607639953
transform 1 0 40462 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_434
timestamp 1607639953
transform 1 0 41014 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_422
timestamp 1607639953
transform 1 0 39910 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_890
timestamp 1607639953
transform 1 0 40370 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_452
timestamp 1607639953
transform 1 0 42670 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_459
timestamp 1607639953
transform 1 0 43314 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_446
timestamp 1607639953
transform 1 0 42118 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_881
timestamp 1607639953
transform 1 0 43222 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_476
timestamp 1607639953
transform 1 0 44878 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_464
timestamp 1607639953
transform 1 0 43774 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_483
timestamp 1607639953
transform 1 0 45522 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_471
timestamp 1607639953
transform 1 0 44418 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_501
timestamp 1607639953
transform 1 0 47178 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_489
timestamp 1607639953
transform 1 0 46074 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_495
timestamp 1607639953
transform 1 0 46626 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_891
timestamp 1607639953
transform 1 0 45982 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_525
timestamp 1607639953
transform 1 0 49386 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_513
timestamp 1607639953
transform 1 0 48282 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_520
timestamp 1607639953
transform 1 0 48926 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_507
timestamp 1607639953
transform 1 0 47730 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_882
timestamp 1607639953
transform 1 0 48834 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_550
timestamp 1607639953
transform 1 0 51686 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_537
timestamp 1607639953
transform 1 0 50490 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_544
timestamp 1607639953
transform 1 0 51134 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_532
timestamp 1607639953
transform 1 0 50030 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_892
timestamp 1607639953
transform 1 0 51594 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_562
timestamp 1607639953
transform 1 0 52790 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_568
timestamp 1607639953
transform 1 0 53342 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_556
timestamp 1607639953
transform 1 0 52238 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_586
timestamp 1607639953
transform 1 0 54998 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_574
timestamp 1607639953
transform 1 0 53894 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_593
timestamp 1607639953
transform 1 0 55642 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_581
timestamp 1607639953
transform 1 0 54538 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_883
timestamp 1607639953
transform 1 0 54446 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_611
timestamp 1607639953
transform 1 0 57298 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_598
timestamp 1607639953
transform 1 0 56102 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_605
timestamp 1607639953
transform 1 0 56746 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_893
timestamp 1607639953
transform 1 0 57206 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_623
timestamp 1607639953
transform 1 0 58402 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_617
timestamp 1607639953
transform 1 0 57850 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1607639953
transform -1 0 58862 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1607639953
transform -1 0 58862 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1607639953
transform 1 0 2466 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1607639953
transform 1 0 1362 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1607639953
transform 1 0 1086 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_44
timestamp 1607639953
transform 1 0 5134 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_32
timestamp 1607639953
transform 1 0 4030 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_27
timestamp 1607639953
transform 1 0 3570 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_894
timestamp 1607639953
transform 1 0 3938 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_56
timestamp 1607639953
transform 1 0 6238 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_80
timestamp 1607639953
transform 1 0 8446 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_68
timestamp 1607639953
transform 1 0 7342 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_105
timestamp 1607639953
transform 1 0 10746 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_93
timestamp 1607639953
transform 1 0 9642 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_895
timestamp 1607639953
transform 1 0 9550 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_129
timestamp 1607639953
transform 1 0 12954 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_117
timestamp 1607639953
transform 1 0 11850 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_154
timestamp 1607639953
transform 1 0 15254 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1607639953
transform 1 0 14058 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_896
timestamp 1607639953
transform 1 0 15162 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_166
timestamp 1607639953
transform 1 0 16358 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_190
timestamp 1607639953
transform 1 0 18566 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_178
timestamp 1607639953
transform 1 0 17462 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_215
timestamp 1607639953
transform 1 0 20866 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_202
timestamp 1607639953
transform 1 0 19670 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_897
timestamp 1607639953
transform 1 0 20774 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_238
timestamp 1607639953
transform 1 0 22982 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_226
timestamp 1607639953
transform 1 0 21878 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _184_
timestamp 1607639953
transform 1 0 21602 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_262
timestamp 1607639953
transform 1 0 25190 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_250
timestamp 1607639953
transform 1 0 24086 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_276
timestamp 1607639953
transform 1 0 26478 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_274
timestamp 1607639953
transform 1 0 26294 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_898
timestamp 1607639953
transform 1 0 26386 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_300
timestamp 1607639953
transform 1 0 28686 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_288
timestamp 1607639953
transform 1 0 27582 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_324
timestamp 1607639953
transform 1 0 30894 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_312
timestamp 1607639953
transform 1 0 29790 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_349
timestamp 1607639953
transform 1 0 33194 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_337
timestamp 1607639953
transform 1 0 32090 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_899
timestamp 1607639953
transform 1 0 31998 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_373
timestamp 1607639953
transform 1 0 35402 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_361
timestamp 1607639953
transform 1 0 34298 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_391
timestamp 1607639953
transform 1 0 37058 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_68_385
timestamp 1607639953
transform 1 0 36506 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _110_
timestamp 1607639953
transform 1 0 36782 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_410
timestamp 1607639953
transform 1 0 38806 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_398
timestamp 1607639953
transform 1 0 37702 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_900
timestamp 1607639953
transform 1 0 37610 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_440
timestamp 1607639953
transform 1 0 41566 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_434
timestamp 1607639953
transform 1 0 41014 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_422
timestamp 1607639953
transform 1 0 39910 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_459
timestamp 1607639953
transform 1 0 43314 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_456
timestamp 1607639953
transform 1 0 43038 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_444
timestamp 1607639953
transform 1 0 41934 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_901
timestamp 1607639953
transform 1 0 43222 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _084_
timestamp 1607639953
transform 1 0 41658 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_483
timestamp 1607639953
transform 1 0 45522 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_471
timestamp 1607639953
transform 1 0 44418 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_495
timestamp 1607639953
transform 1 0 46626 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_520
timestamp 1607639953
transform 1 0 48926 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_507
timestamp 1607639953
transform 1 0 47730 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_902
timestamp 1607639953
transform 1 0 48834 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_544
timestamp 1607639953
transform 1 0 51134 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_532
timestamp 1607639953
transform 1 0 50030 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_568
timestamp 1607639953
transform 1 0 53342 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_556
timestamp 1607639953
transform 1 0 52238 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_593
timestamp 1607639953
transform 1 0 55642 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_581
timestamp 1607639953
transform 1 0 54538 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_903
timestamp 1607639953
transform 1 0 54446 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_611
timestamp 1607639953
transform 1 0 57298 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_599
timestamp 1607639953
transform 1 0 56194 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _144_
timestamp 1607639953
transform 1 0 55918 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_623
timestamp 1607639953
transform 1 0 58402 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1607639953
transform -1 0 58862 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1607639953
transform 1 0 2466 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1607639953
transform 1 0 1362 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1607639953
transform 1 0 1086 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_43
timestamp 1607639953
transform 1 0 5042 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_39
timestamp 1607639953
transform 1 0 4674 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1607639953
transform 1 0 3570 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _189_
timestamp 1607639953
transform 1 0 4766 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_62
timestamp 1607639953
transform 1 0 6790 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_55
timestamp 1607639953
transform 1 0 6146 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_904
timestamp 1607639953
transform 1 0 6698 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_86
timestamp 1607639953
transform 1 0 8998 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_74
timestamp 1607639953
transform 1 0 7894 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_110
timestamp 1607639953
transform 1 0 11206 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_98
timestamp 1607639953
transform 1 0 10102 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_123
timestamp 1607639953
transform 1 0 12402 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_905
timestamp 1607639953
transform 1 0 12310 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_148
timestamp 1607639953
transform 1 0 14702 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_143
timestamp 1607639953
transform 1 0 14242 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_135
timestamp 1607639953
transform 1 0 13506 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _108_
timestamp 1607639953
transform 1 0 14426 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_172
timestamp 1607639953
transform 1 0 16910 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_160
timestamp 1607639953
transform 1 0 15806 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_196
timestamp 1607639953
transform 1 0 19118 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_184
timestamp 1607639953
transform 1 0 18014 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_180
timestamp 1607639953
transform 1 0 17646 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_906
timestamp 1607639953
transform 1 0 17922 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_220
timestamp 1607639953
transform 1 0 21326 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_208
timestamp 1607639953
transform 1 0 20222 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_232
timestamp 1607639953
transform 1 0 22430 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_257
timestamp 1607639953
transform 1 0 24730 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_245
timestamp 1607639953
transform 1 0 23626 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_907
timestamp 1607639953
transform 1 0 23534 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1607639953
transform 1 0 26938 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_269
timestamp 1607639953
transform 1 0 25834 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_306
timestamp 1607639953
transform 1 0 29238 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1607639953
transform 1 0 28042 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_908
timestamp 1607639953
transform 1 0 29146 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_330
timestamp 1607639953
transform 1 0 31446 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_318
timestamp 1607639953
transform 1 0 30342 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_342
timestamp 1607639953
transform 1 0 32550 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_367
timestamp 1607639953
transform 1 0 34850 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_354
timestamp 1607639953
transform 1 0 33654 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_909
timestamp 1607639953
transform 1 0 34758 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_391
timestamp 1607639953
transform 1 0 37058 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_379
timestamp 1607639953
transform 1 0 35954 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_415
timestamp 1607639953
transform 1 0 39266 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_403
timestamp 1607639953
transform 1 0 38162 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_440
timestamp 1607639953
transform 1 0 41566 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_428
timestamp 1607639953
transform 1 0 40462 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_910
timestamp 1607639953
transform 1 0 40370 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_452
timestamp 1607639953
transform 1 0 42670 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_476
timestamp 1607639953
transform 1 0 44878 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_464
timestamp 1607639953
transform 1 0 43774 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_501
timestamp 1607639953
transform 1 0 47178 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_489
timestamp 1607639953
transform 1 0 46074 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_911
timestamp 1607639953
transform 1 0 45982 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_525
timestamp 1607639953
transform 1 0 49386 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_513
timestamp 1607639953
transform 1 0 48282 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_550
timestamp 1607639953
transform 1 0 51686 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_537
timestamp 1607639953
transform 1 0 50490 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_912
timestamp 1607639953
transform 1 0 51594 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_562
timestamp 1607639953
transform 1 0 52790 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_586
timestamp 1607639953
transform 1 0 54998 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_574
timestamp 1607639953
transform 1 0 53894 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_615
timestamp 1607639953
transform 1 0 57666 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_611
timestamp 1607639953
transform 1 0 57298 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_598
timestamp 1607639953
transform 1 0 56102 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_913
timestamp 1607639953
transform 1 0 57206 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _089_
timestamp 1607639953
transform 1 0 57390 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_623
timestamp 1607639953
transform 1 0 58402 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1607639953
transform -1 0 58862 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1607639953
transform 1 0 2466 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1607639953
transform 1 0 1362 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1607639953
transform 1 0 1086 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_44
timestamp 1607639953
transform 1 0 5134 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_32
timestamp 1607639953
transform 1 0 4030 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_27
timestamp 1607639953
transform 1 0 3570 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_914
timestamp 1607639953
transform 1 0 3938 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_59
timestamp 1607639953
transform 1 0 6514 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _099_
timestamp 1607639953
transform 1 0 6238 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_83
timestamp 1607639953
transform 1 0 8722 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_71
timestamp 1607639953
transform 1 0 7618 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_105
timestamp 1607639953
transform 1 0 10746 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_93
timestamp 1607639953
transform 1 0 9642 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_91
timestamp 1607639953
transform 1 0 9458 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_915
timestamp 1607639953
transform 1 0 9550 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_129
timestamp 1607639953
transform 1 0 12954 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_117
timestamp 1607639953
transform 1 0 11850 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_154
timestamp 1607639953
transform 1 0 15254 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1607639953
transform 1 0 14058 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_916
timestamp 1607639953
transform 1 0 15162 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_166
timestamp 1607639953
transform 1 0 16358 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_190
timestamp 1607639953
transform 1 0 18566 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_178
timestamp 1607639953
transform 1 0 17462 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_215
timestamp 1607639953
transform 1 0 20866 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_202
timestamp 1607639953
transform 1 0 19670 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_917
timestamp 1607639953
transform 1 0 20774 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_239
timestamp 1607639953
transform 1 0 23074 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_227
timestamp 1607639953
transform 1 0 21970 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_263
timestamp 1607639953
transform 1 0 25282 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_251
timestamp 1607639953
transform 1 0 24178 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_276
timestamp 1607639953
transform 1 0 26478 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_918
timestamp 1607639953
transform 1 0 26386 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_300
timestamp 1607639953
transform 1 0 28686 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_288
timestamp 1607639953
transform 1 0 27582 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_324
timestamp 1607639953
transform 1 0 30894 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_312
timestamp 1607639953
transform 1 0 29790 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_349
timestamp 1607639953
transform 1 0 33194 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_337
timestamp 1607639953
transform 1 0 32090 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_919
timestamp 1607639953
transform 1 0 31998 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_373
timestamp 1607639953
transform 1 0 35402 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_361
timestamp 1607639953
transform 1 0 34298 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_385
timestamp 1607639953
transform 1 0 36506 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_410
timestamp 1607639953
transform 1 0 38806 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_398
timestamp 1607639953
transform 1 0 37702 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_920
timestamp 1607639953
transform 1 0 37610 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_434
timestamp 1607639953
transform 1 0 41014 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_422
timestamp 1607639953
transform 1 0 39910 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_459
timestamp 1607639953
transform 1 0 43314 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_446
timestamp 1607639953
transform 1 0 42118 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_921
timestamp 1607639953
transform 1 0 43222 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_483
timestamp 1607639953
transform 1 0 45522 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_471
timestamp 1607639953
transform 1 0 44418 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_495
timestamp 1607639953
transform 1 0 46626 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_520
timestamp 1607639953
transform 1 0 48926 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_507
timestamp 1607639953
transform 1 0 47730 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_922
timestamp 1607639953
transform 1 0 48834 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_544
timestamp 1607639953
transform 1 0 51134 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_532
timestamp 1607639953
transform 1 0 50030 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_568
timestamp 1607639953
transform 1 0 53342 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_556
timestamp 1607639953
transform 1 0 52238 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_593
timestamp 1607639953
transform 1 0 55642 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_581
timestamp 1607639953
transform 1 0 54538 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_923
timestamp 1607639953
transform 1 0 54446 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _145_
timestamp 1607639953
transform 1 0 55734 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_609
timestamp 1607639953
transform 1 0 57114 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_597
timestamp 1607639953
transform 1 0 56010 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_621
timestamp 1607639953
transform 1 0 58218 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1607639953
transform -1 0 58862 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1607639953
transform 1 0 2466 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1607639953
transform 1 0 1362 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1607639953
transform 1 0 1086 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1607639953
transform 1 0 4674 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1607639953
transform 1 0 3570 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_62
timestamp 1607639953
transform 1 0 6790 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_71_59
timestamp 1607639953
transform 1 0 6514 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_51
timestamp 1607639953
transform 1 0 5778 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_924
timestamp 1607639953
transform 1 0 6698 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_83
timestamp 1607639953
transform 1 0 8722 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_71
timestamp 1607639953
transform 1 0 7618 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _086_
timestamp 1607639953
transform 1 0 7342 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_110
timestamp 1607639953
transform 1 0 11206 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_95
timestamp 1607639953
transform 1 0 9826 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _101_
timestamp 1607639953
transform 1 0 10930 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_123
timestamp 1607639953
transform 1 0 12402 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_925
timestamp 1607639953
transform 1 0 12310 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_147
timestamp 1607639953
transform 1 0 14610 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_135
timestamp 1607639953
transform 1 0 13506 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_171
timestamp 1607639953
transform 1 0 16818 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_159
timestamp 1607639953
transform 1 0 15714 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_196
timestamp 1607639953
transform 1 0 19118 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_184
timestamp 1607639953
transform 1 0 18014 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_926
timestamp 1607639953
transform 1 0 17922 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_218
timestamp 1607639953
transform 1 0 21142 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_206
timestamp 1607639953
transform 1 0 20038 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_202
timestamp 1607639953
transform 1 0 19670 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1607639953
transform 1 0 19762 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_242
timestamp 1607639953
transform 1 0 23350 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_230
timestamp 1607639953
transform 1 0 22246 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_257
timestamp 1607639953
transform 1 0 24730 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_245
timestamp 1607639953
transform 1 0 23626 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_927
timestamp 1607639953
transform 1 0 23534 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1607639953
transform 1 0 26938 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_269
timestamp 1607639953
transform 1 0 25834 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_306
timestamp 1607639953
transform 1 0 29238 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1607639953
transform 1 0 28042 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_928
timestamp 1607639953
transform 1 0 29146 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_330
timestamp 1607639953
transform 1 0 31446 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_318
timestamp 1607639953
transform 1 0 30342 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_342
timestamp 1607639953
transform 1 0 32550 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_367
timestamp 1607639953
transform 1 0 34850 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_354
timestamp 1607639953
transform 1 0 33654 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_929
timestamp 1607639953
transform 1 0 34758 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_391
timestamp 1607639953
transform 1 0 37058 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_379
timestamp 1607639953
transform 1 0 35954 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_415
timestamp 1607639953
transform 1 0 39266 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_403
timestamp 1607639953
transform 1 0 38162 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_440
timestamp 1607639953
transform 1 0 41566 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_428
timestamp 1607639953
transform 1 0 40462 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_930
timestamp 1607639953
transform 1 0 40370 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_452
timestamp 1607639953
transform 1 0 42670 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_476
timestamp 1607639953
transform 1 0 44878 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_464
timestamp 1607639953
transform 1 0 43774 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_501
timestamp 1607639953
transform 1 0 47178 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_489
timestamp 1607639953
transform 1 0 46074 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_931
timestamp 1607639953
transform 1 0 45982 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_525
timestamp 1607639953
transform 1 0 49386 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_513
timestamp 1607639953
transform 1 0 48282 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_550
timestamp 1607639953
transform 1 0 51686 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_537
timestamp 1607639953
transform 1 0 50490 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_932
timestamp 1607639953
transform 1 0 51594 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_562
timestamp 1607639953
transform 1 0 52790 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_586
timestamp 1607639953
transform 1 0 54998 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_574
timestamp 1607639953
transform 1 0 53894 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_611
timestamp 1607639953
transform 1 0 57298 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_598
timestamp 1607639953
transform 1 0 56102 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_933
timestamp 1607639953
transform 1 0 57206 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_623
timestamp 1607639953
transform 1 0 58402 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1607639953
transform -1 0 58862 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1607639953
transform 1 0 2466 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1607639953
transform 1 0 1362 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1607639953
transform 1 0 2466 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1607639953
transform 1 0 1362 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1607639953
transform 1 0 1086 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1607639953
transform 1 0 1086 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1607639953
transform 1 0 4674 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1607639953
transform 1 0 3570 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_44
timestamp 1607639953
transform 1 0 5134 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_32
timestamp 1607639953
transform 1 0 4030 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_27
timestamp 1607639953
transform 1 0 3570 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_934
timestamp 1607639953
transform 1 0 3938 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_62
timestamp 1607639953
transform 1 0 6790 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_59
timestamp 1607639953
transform 1 0 6514 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_51
timestamp 1607639953
transform 1 0 5778 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_56
timestamp 1607639953
transform 1 0 6238 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_944
timestamp 1607639953
transform 1 0 6698 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_86
timestamp 1607639953
transform 1 0 8998 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_74
timestamp 1607639953
transform 1 0 7894 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_80
timestamp 1607639953
transform 1 0 8446 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_68
timestamp 1607639953
transform 1 0 7342 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_99
timestamp 1607639953
transform 1 0 10194 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_94
timestamp 1607639953
transform 1 0 9734 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_105
timestamp 1607639953
transform 1 0 10746 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_93
timestamp 1607639953
transform 1 0 9642 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_935
timestamp 1607639953
transform 1 0 9550 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _018_
timestamp 1607639953
transform 1 0 9918 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_123
timestamp 1607639953
transform 1 0 12402 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_119
timestamp 1607639953
transform 1 0 12034 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_111
timestamp 1607639953
transform 1 0 11298 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_129
timestamp 1607639953
transform 1 0 12954 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_117
timestamp 1607639953
transform 1 0 11850 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_945
timestamp 1607639953
transform 1 0 12310 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_147
timestamp 1607639953
transform 1 0 14610 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_135
timestamp 1607639953
transform 1 0 13506 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_154
timestamp 1607639953
transform 1 0 15254 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1607639953
transform 1 0 14058 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_936
timestamp 1607639953
transform 1 0 15162 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_171
timestamp 1607639953
transform 1 0 16818 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_159
timestamp 1607639953
transform 1 0 15714 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_166
timestamp 1607639953
transform 1 0 16358 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_196
timestamp 1607639953
transform 1 0 19118 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_184
timestamp 1607639953
transform 1 0 18014 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_190
timestamp 1607639953
transform 1 0 18566 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_178
timestamp 1607639953
transform 1 0 17462 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_946
timestamp 1607639953
transform 1 0 17922 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_220
timestamp 1607639953
transform 1 0 21326 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_208
timestamp 1607639953
transform 1 0 20222 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_215
timestamp 1607639953
transform 1 0 20866 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_202
timestamp 1607639953
transform 1 0 19670 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_937
timestamp 1607639953
transform 1 0 20774 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_232
timestamp 1607639953
transform 1 0 22430 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_239
timestamp 1607639953
transform 1 0 23074 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_227
timestamp 1607639953
transform 1 0 21970 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_257
timestamp 1607639953
transform 1 0 24730 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_245
timestamp 1607639953
transform 1 0 23626 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_263
timestamp 1607639953
transform 1 0 25282 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_251
timestamp 1607639953
transform 1 0 24178 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_947
timestamp 1607639953
transform 1 0 23534 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1607639953
transform 1 0 26938 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_269
timestamp 1607639953
transform 1 0 25834 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_276
timestamp 1607639953
transform 1 0 26478 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_938
timestamp 1607639953
transform 1 0 26386 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_306
timestamp 1607639953
transform 1 0 29238 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1607639953
transform 1 0 28042 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_300
timestamp 1607639953
transform 1 0 28686 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_288
timestamp 1607639953
transform 1 0 27582 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_948
timestamp 1607639953
transform 1 0 29146 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_330
timestamp 1607639953
transform 1 0 31446 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_318
timestamp 1607639953
transform 1 0 30342 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_324
timestamp 1607639953
transform 1 0 30894 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_312
timestamp 1607639953
transform 1 0 29790 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_342
timestamp 1607639953
transform 1 0 32550 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_349
timestamp 1607639953
transform 1 0 33194 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_337
timestamp 1607639953
transform 1 0 32090 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_939
timestamp 1607639953
transform 1 0 31998 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_367
timestamp 1607639953
transform 1 0 34850 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_354
timestamp 1607639953
transform 1 0 33654 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_373
timestamp 1607639953
transform 1 0 35402 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_361
timestamp 1607639953
transform 1 0 34298 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_949
timestamp 1607639953
transform 1 0 34758 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1607639953
transform 1 0 37242 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_381
timestamp 1607639953
transform 1 0 36138 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_375
timestamp 1607639953
transform 1 0 35586 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_385
timestamp 1607639953
transform 1 0 36506 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _205_
timestamp 1607639953
transform 1 0 35862 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_417
timestamp 1607639953
transform 1 0 39450 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1607639953
transform 1 0 38346 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_410
timestamp 1607639953
transform 1 0 38806 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_398
timestamp 1607639953
transform 1 0 37702 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_940
timestamp 1607639953
transform 1 0 37610 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_440
timestamp 1607639953
transform 1 0 41566 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_428
timestamp 1607639953
transform 1 0 40462 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_425
timestamp 1607639953
transform 1 0 40186 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_434
timestamp 1607639953
transform 1 0 41014 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_422
timestamp 1607639953
transform 1 0 39910 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_950
timestamp 1607639953
transform 1 0 40370 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_452
timestamp 1607639953
transform 1 0 42670 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_459
timestamp 1607639953
transform 1 0 43314 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_446
timestamp 1607639953
transform 1 0 42118 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_941
timestamp 1607639953
transform 1 0 43222 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_476
timestamp 1607639953
transform 1 0 44878 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_464
timestamp 1607639953
transform 1 0 43774 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_483
timestamp 1607639953
transform 1 0 45522 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_471
timestamp 1607639953
transform 1 0 44418 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_501
timestamp 1607639953
transform 1 0 47178 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_489
timestamp 1607639953
transform 1 0 46074 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_495
timestamp 1607639953
transform 1 0 46626 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_951
timestamp 1607639953
transform 1 0 45982 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_525
timestamp 1607639953
transform 1 0 49386 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_513
timestamp 1607639953
transform 1 0 48282 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_520
timestamp 1607639953
transform 1 0 48926 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_507
timestamp 1607639953
transform 1 0 47730 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_942
timestamp 1607639953
transform 1 0 48834 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_550
timestamp 1607639953
transform 1 0 51686 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_537
timestamp 1607639953
transform 1 0 50490 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_544
timestamp 1607639953
transform 1 0 51134 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_532
timestamp 1607639953
transform 1 0 50030 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_952
timestamp 1607639953
transform 1 0 51594 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_562
timestamp 1607639953
transform 1 0 52790 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_568
timestamp 1607639953
transform 1 0 53342 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_556
timestamp 1607639953
transform 1 0 52238 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_586
timestamp 1607639953
transform 1 0 54998 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_574
timestamp 1607639953
transform 1 0 53894 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_593
timestamp 1607639953
transform 1 0 55642 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_581
timestamp 1607639953
transform 1 0 54538 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_943
timestamp 1607639953
transform 1 0 54446 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_611
timestamp 1607639953
transform 1 0 57298 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_598
timestamp 1607639953
transform 1 0 56102 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_605
timestamp 1607639953
transform 1 0 56746 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_953
timestamp 1607639953
transform 1 0 57206 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_623
timestamp 1607639953
transform 1 0 58402 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_617
timestamp 1607639953
transform 1 0 57850 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1607639953
transform -1 0 58862 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1607639953
transform -1 0 58862 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1607639953
transform 1 0 2466 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1607639953
transform 1 0 1362 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1607639953
transform 1 0 1086 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_44
timestamp 1607639953
transform 1 0 5134 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_32
timestamp 1607639953
transform 1 0 4030 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_27
timestamp 1607639953
transform 1 0 3570 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_954
timestamp 1607639953
transform 1 0 3938 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_56
timestamp 1607639953
transform 1 0 6238 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_80
timestamp 1607639953
transform 1 0 8446 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_68
timestamp 1607639953
transform 1 0 7342 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_105
timestamp 1607639953
transform 1 0 10746 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_93
timestamp 1607639953
transform 1 0 9642 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_955
timestamp 1607639953
transform 1 0 9550 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_129
timestamp 1607639953
transform 1 0 12954 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_117
timestamp 1607639953
transform 1 0 11850 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_154
timestamp 1607639953
transform 1 0 15254 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1607639953
transform 1 0 14058 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_956
timestamp 1607639953
transform 1 0 15162 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_166
timestamp 1607639953
transform 1 0 16358 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_190
timestamp 1607639953
transform 1 0 18566 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_178
timestamp 1607639953
transform 1 0 17462 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_215
timestamp 1607639953
transform 1 0 20866 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_202
timestamp 1607639953
transform 1 0 19670 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_957
timestamp 1607639953
transform 1 0 20774 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_239
timestamp 1607639953
transform 1 0 23074 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_227
timestamp 1607639953
transform 1 0 21970 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_263
timestamp 1607639953
transform 1 0 25282 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_251
timestamp 1607639953
transform 1 0 24178 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_276
timestamp 1607639953
transform 1 0 26478 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_958
timestamp 1607639953
transform 1 0 26386 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_300
timestamp 1607639953
transform 1 0 28686 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_288
timestamp 1607639953
transform 1 0 27582 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_324
timestamp 1607639953
transform 1 0 30894 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_312
timestamp 1607639953
transform 1 0 29790 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_349
timestamp 1607639953
transform 1 0 33194 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_337
timestamp 1607639953
transform 1 0 32090 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_959
timestamp 1607639953
transform 1 0 31998 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_373
timestamp 1607639953
transform 1 0 35402 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_361
timestamp 1607639953
transform 1 0 34298 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_385
timestamp 1607639953
transform 1 0 36506 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_410
timestamp 1607639953
transform 1 0 38806 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_398
timestamp 1607639953
transform 1 0 37702 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_960
timestamp 1607639953
transform 1 0 37610 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_434
timestamp 1607639953
transform 1 0 41014 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_422
timestamp 1607639953
transform 1 0 39910 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_459
timestamp 1607639953
transform 1 0 43314 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_446
timestamp 1607639953
transform 1 0 42118 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_961
timestamp 1607639953
transform 1 0 43222 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_483
timestamp 1607639953
transform 1 0 45522 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_471
timestamp 1607639953
transform 1 0 44418 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_495
timestamp 1607639953
transform 1 0 46626 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_520
timestamp 1607639953
transform 1 0 48926 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_507
timestamp 1607639953
transform 1 0 47730 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_962
timestamp 1607639953
transform 1 0 48834 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_544
timestamp 1607639953
transform 1 0 51134 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_532
timestamp 1607639953
transform 1 0 50030 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_568
timestamp 1607639953
transform 1 0 53342 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_556
timestamp 1607639953
transform 1 0 52238 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_593
timestamp 1607639953
transform 1 0 55642 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_581
timestamp 1607639953
transform 1 0 54538 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_963
timestamp 1607639953
transform 1 0 54446 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_605
timestamp 1607639953
transform 1 0 56746 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_617
timestamp 1607639953
transform 1 0 57850 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1607639953
transform -1 0 58862 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_18
timestamp 1607639953
transform 1 0 2742 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_6
timestamp 1607639953
transform 1 0 1638 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1607639953
transform 1 0 1086 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _003_
timestamp 1607639953
transform 1 0 1362 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_42
timestamp 1607639953
transform 1 0 4950 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_30
timestamp 1607639953
transform 1 0 3846 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_62
timestamp 1607639953
transform 1 0 6790 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_60
timestamp 1607639953
transform 1 0 6606 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_54
timestamp 1607639953
transform 1 0 6054 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_964
timestamp 1607639953
transform 1 0 6698 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_86
timestamp 1607639953
transform 1 0 8998 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_74
timestamp 1607639953
transform 1 0 7894 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_99
timestamp 1607639953
transform 1 0 10194 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_94
timestamp 1607639953
transform 1 0 9734 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _013_
timestamp 1607639953
transform 1 0 9918 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_123
timestamp 1607639953
transform 1 0 12402 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_119
timestamp 1607639953
transform 1 0 12034 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_111
timestamp 1607639953
transform 1 0 11298 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_965
timestamp 1607639953
transform 1 0 12310 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_152
timestamp 1607639953
transform 1 0 15070 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_147
timestamp 1607639953
transform 1 0 14610 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_135
timestamp 1607639953
transform 1 0 13506 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1607639953
transform 1 0 14794 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_176
timestamp 1607639953
transform 1 0 17278 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_164
timestamp 1607639953
transform 1 0 16174 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_196
timestamp 1607639953
transform 1 0 19118 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_184
timestamp 1607639953
transform 1 0 18014 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_182
timestamp 1607639953
transform 1 0 17830 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_966
timestamp 1607639953
transform 1 0 17922 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_220
timestamp 1607639953
transform 1 0 21326 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_208
timestamp 1607639953
transform 1 0 20222 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_232
timestamp 1607639953
transform 1 0 22430 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_257
timestamp 1607639953
transform 1 0 24730 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_245
timestamp 1607639953
transform 1 0 23626 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_967
timestamp 1607639953
transform 1 0 23534 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1607639953
transform 1 0 26938 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_269
timestamp 1607639953
transform 1 0 25834 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_306
timestamp 1607639953
transform 1 0 29238 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1607639953
transform 1 0 28042 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_968
timestamp 1607639953
transform 1 0 29146 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_330
timestamp 1607639953
transform 1 0 31446 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_318
timestamp 1607639953
transform 1 0 30342 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_342
timestamp 1607639953
transform 1 0 32550 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_367
timestamp 1607639953
transform 1 0 34850 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_354
timestamp 1607639953
transform 1 0 33654 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_969
timestamp 1607639953
transform 1 0 34758 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_391
timestamp 1607639953
transform 1 0 37058 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_379
timestamp 1607639953
transform 1 0 35954 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_415
timestamp 1607639953
transform 1 0 39266 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_403
timestamp 1607639953
transform 1 0 38162 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_440
timestamp 1607639953
transform 1 0 41566 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_428
timestamp 1607639953
transform 1 0 40462 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_970
timestamp 1607639953
transform 1 0 40370 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_452
timestamp 1607639953
transform 1 0 42670 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_476
timestamp 1607639953
transform 1 0 44878 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_464
timestamp 1607639953
transform 1 0 43774 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_501
timestamp 1607639953
transform 1 0 47178 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_489
timestamp 1607639953
transform 1 0 46074 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_971
timestamp 1607639953
transform 1 0 45982 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_525
timestamp 1607639953
transform 1 0 49386 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_513
timestamp 1607639953
transform 1 0 48282 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_550
timestamp 1607639953
transform 1 0 51686 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_537
timestamp 1607639953
transform 1 0 50490 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_972
timestamp 1607639953
transform 1 0 51594 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_562
timestamp 1607639953
transform 1 0 52790 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_586
timestamp 1607639953
transform 1 0 54998 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_574
timestamp 1607639953
transform 1 0 53894 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_611
timestamp 1607639953
transform 1 0 57298 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_598
timestamp 1607639953
transform 1 0 56102 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_973
timestamp 1607639953
transform 1 0 57206 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_623
timestamp 1607639953
transform 1 0 58402 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1607639953
transform -1 0 58862 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1607639953
transform 1 0 2466 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1607639953
transform 1 0 1362 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1607639953
transform 1 0 1086 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_44
timestamp 1607639953
transform 1 0 5134 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_32
timestamp 1607639953
transform 1 0 4030 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_27
timestamp 1607639953
transform 1 0 3570 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_974
timestamp 1607639953
transform 1 0 3938 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_62
timestamp 1607639953
transform 1 0 6790 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_56
timestamp 1607639953
transform 1 0 6238 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _074_
timestamp 1607639953
transform 1 0 6514 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_76_86
timestamp 1607639953
transform 1 0 8998 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_74
timestamp 1607639953
transform 1 0 7894 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_105
timestamp 1607639953
transform 1 0 10746 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_93
timestamp 1607639953
transform 1 0 9642 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_975
timestamp 1607639953
transform 1 0 9550 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_129
timestamp 1607639953
transform 1 0 12954 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_117
timestamp 1607639953
transform 1 0 11850 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_154
timestamp 1607639953
transform 1 0 15254 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1607639953
transform 1 0 14058 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_976
timestamp 1607639953
transform 1 0 15162 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_166
timestamp 1607639953
transform 1 0 16358 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_190
timestamp 1607639953
transform 1 0 18566 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_178
timestamp 1607639953
transform 1 0 17462 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_215
timestamp 1607639953
transform 1 0 20866 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_202
timestamp 1607639953
transform 1 0 19670 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_977
timestamp 1607639953
transform 1 0 20774 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_239
timestamp 1607639953
transform 1 0 23074 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_227
timestamp 1607639953
transform 1 0 21970 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_263
timestamp 1607639953
transform 1 0 25282 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_251
timestamp 1607639953
transform 1 0 24178 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_276
timestamp 1607639953
transform 1 0 26478 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_978
timestamp 1607639953
transform 1 0 26386 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_300
timestamp 1607639953
transform 1 0 28686 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_288
timestamp 1607639953
transform 1 0 27582 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_324
timestamp 1607639953
transform 1 0 30894 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_312
timestamp 1607639953
transform 1 0 29790 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_349
timestamp 1607639953
transform 1 0 33194 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_337
timestamp 1607639953
transform 1 0 32090 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_979
timestamp 1607639953
transform 1 0 31998 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_373
timestamp 1607639953
transform 1 0 35402 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_361
timestamp 1607639953
transform 1 0 34298 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_396
timestamp 1607639953
transform 1 0 37518 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_385
timestamp 1607639953
transform 1 0 36506 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _136_
timestamp 1607639953
transform 1 0 37242 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_410
timestamp 1607639953
transform 1 0 38806 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_398
timestamp 1607639953
transform 1 0 37702 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_980
timestamp 1607639953
transform 1 0 37610 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_434
timestamp 1607639953
transform 1 0 41014 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_422
timestamp 1607639953
transform 1 0 39910 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_459
timestamp 1607639953
transform 1 0 43314 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_446
timestamp 1607639953
transform 1 0 42118 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_981
timestamp 1607639953
transform 1 0 43222 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_479
timestamp 1607639953
transform 1 0 45154 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1607639953
transform 1 0 44786 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_471
timestamp 1607639953
transform 1 0 44418 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _012_
timestamp 1607639953
transform 1 0 44878 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_503
timestamp 1607639953
transform 1 0 47362 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_491
timestamp 1607639953
transform 1 0 46258 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_520
timestamp 1607639953
transform 1 0 48926 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_515
timestamp 1607639953
transform 1 0 48466 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_982
timestamp 1607639953
transform 1 0 48834 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_550
timestamp 1607639953
transform 1 0 51686 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_544
timestamp 1607639953
transform 1 0 51134 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_532
timestamp 1607639953
transform 1 0 50030 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_565
timestamp 1607639953
transform 1 0 53066 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_554
timestamp 1607639953
transform 1 0 52054 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _071_
timestamp 1607639953
transform 1 0 52790 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _025_
timestamp 1607639953
transform 1 0 51778 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_593
timestamp 1607639953
transform 1 0 55642 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_581
timestamp 1607639953
transform 1 0 54538 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_577
timestamp 1607639953
transform 1 0 54170 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_983
timestamp 1607639953
transform 1 0 54446 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_605
timestamp 1607639953
transform 1 0 56746 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_617
timestamp 1607639953
transform 1 0 57850 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1607639953
transform -1 0 58862 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1607639953
transform 1 0 2466 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1607639953
transform 1 0 1362 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1607639953
transform 1 0 1086 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1607639953
transform 1 0 4674 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1607639953
transform 1 0 3570 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_62
timestamp 1607639953
transform 1 0 6790 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_59
timestamp 1607639953
transform 1 0 6514 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_51
timestamp 1607639953
transform 1 0 5778 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_984
timestamp 1607639953
transform 1 0 6698 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_86
timestamp 1607639953
transform 1 0 8998 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_74
timestamp 1607639953
transform 1 0 7894 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_110
timestamp 1607639953
transform 1 0 11206 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_98
timestamp 1607639953
transform 1 0 10102 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_123
timestamp 1607639953
transform 1 0 12402 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_985
timestamp 1607639953
transform 1 0 12310 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_151
timestamp 1607639953
transform 1 0 14978 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_139
timestamp 1607639953
transform 1 0 13874 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_135
timestamp 1607639953
transform 1 0 13506 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _090_
timestamp 1607639953
transform 1 0 13598 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_175
timestamp 1607639953
transform 1 0 17186 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_163
timestamp 1607639953
transform 1 0 16082 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_196
timestamp 1607639953
transform 1 0 19118 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_184
timestamp 1607639953
transform 1 0 18014 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_986
timestamp 1607639953
transform 1 0 17922 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_220
timestamp 1607639953
transform 1 0 21326 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_208
timestamp 1607639953
transform 1 0 20222 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_232
timestamp 1607639953
transform 1 0 22430 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_257
timestamp 1607639953
transform 1 0 24730 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_245
timestamp 1607639953
transform 1 0 23626 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_987
timestamp 1607639953
transform 1 0 23534 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1607639953
transform 1 0 26938 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_269
timestamp 1607639953
transform 1 0 25834 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_306
timestamp 1607639953
transform 1 0 29238 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1607639953
transform 1 0 28042 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_988
timestamp 1607639953
transform 1 0 29146 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_327
timestamp 1607639953
transform 1 0 31170 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_315
timestamp 1607639953
transform 1 0 30066 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _111_
timestamp 1607639953
transform 1 0 29790 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_351
timestamp 1607639953
transform 1 0 33378 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_339
timestamp 1607639953
transform 1 0 32274 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_367
timestamp 1607639953
transform 1 0 34850 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_363
timestamp 1607639953
transform 1 0 34482 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_989
timestamp 1607639953
transform 1 0 34758 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_387
timestamp 1607639953
transform 1 0 36690 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_383
timestamp 1607639953
transform 1 0 36322 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_379
timestamp 1607639953
transform 1 0 35954 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _116_
timestamp 1607639953
transform 1 0 36414 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_416
timestamp 1607639953
transform 1 0 39358 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_404
timestamp 1607639953
transform 1 0 38254 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_399
timestamp 1607639953
transform 1 0 37794 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _126_
timestamp 1607639953
transform 1 0 37978 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_440
timestamp 1607639953
transform 1 0 41566 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_428
timestamp 1607639953
transform 1 0 40462 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_424
timestamp 1607639953
transform 1 0 40094 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_990
timestamp 1607639953
transform 1 0 40370 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_451
timestamp 1607639953
transform 1 0 42578 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _183_
timestamp 1607639953
transform 1 0 42302 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_475
timestamp 1607639953
transform 1 0 44786 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_463
timestamp 1607639953
transform 1 0 43682 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_501
timestamp 1607639953
transform 1 0 47178 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_489
timestamp 1607639953
transform 1 0 46074 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_487
timestamp 1607639953
transform 1 0 45890 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_991
timestamp 1607639953
transform 1 0 45982 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_525
timestamp 1607639953
transform 1 0 49386 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_513
timestamp 1607639953
transform 1 0 48282 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_550
timestamp 1607639953
transform 1 0 51686 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_537
timestamp 1607639953
transform 1 0 50490 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_992
timestamp 1607639953
transform 1 0 51594 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_562
timestamp 1607639953
transform 1 0 52790 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_586
timestamp 1607639953
transform 1 0 54998 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_574
timestamp 1607639953
transform 1 0 53894 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_611
timestamp 1607639953
transform 1 0 57298 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_598
timestamp 1607639953
transform 1 0 56102 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_993
timestamp 1607639953
transform 1 0 57206 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_623
timestamp 1607639953
transform 1 0 58402 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1607639953
transform -1 0 58862 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1607639953
transform 1 0 2466 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1607639953
transform 1 0 1362 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1607639953
transform 1 0 1086 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_44
timestamp 1607639953
transform 1 0 5134 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_32
timestamp 1607639953
transform 1 0 4030 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_27
timestamp 1607639953
transform 1 0 3570 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_994
timestamp 1607639953
transform 1 0 3938 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_56
timestamp 1607639953
transform 1 0 6238 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_80
timestamp 1607639953
transform 1 0 8446 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_68
timestamp 1607639953
transform 1 0 7342 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_105
timestamp 1607639953
transform 1 0 10746 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_93
timestamp 1607639953
transform 1 0 9642 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_995
timestamp 1607639953
transform 1 0 9550 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_129
timestamp 1607639953
transform 1 0 12954 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_117
timestamp 1607639953
transform 1 0 11850 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_154
timestamp 1607639953
transform 1 0 15254 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1607639953
transform 1 0 14058 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_996
timestamp 1607639953
transform 1 0 15162 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_166
timestamp 1607639953
transform 1 0 16358 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_190
timestamp 1607639953
transform 1 0 18566 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_178
timestamp 1607639953
transform 1 0 17462 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_215
timestamp 1607639953
transform 1 0 20866 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_202
timestamp 1607639953
transform 1 0 19670 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_997
timestamp 1607639953
transform 1 0 20774 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_239
timestamp 1607639953
transform 1 0 23074 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_227
timestamp 1607639953
transform 1 0 21970 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_263
timestamp 1607639953
transform 1 0 25282 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_251
timestamp 1607639953
transform 1 0 24178 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_276
timestamp 1607639953
transform 1 0 26478 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_998
timestamp 1607639953
transform 1 0 26386 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_300
timestamp 1607639953
transform 1 0 28686 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_288
timestamp 1607639953
transform 1 0 27582 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_324
timestamp 1607639953
transform 1 0 30894 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_312
timestamp 1607639953
transform 1 0 29790 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_349
timestamp 1607639953
transform 1 0 33194 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_337
timestamp 1607639953
transform 1 0 32090 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_999
timestamp 1607639953
transform 1 0 31998 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_373
timestamp 1607639953
transform 1 0 35402 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_361
timestamp 1607639953
transform 1 0 34298 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_396
timestamp 1607639953
transform 1 0 37518 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_390
timestamp 1607639953
transform 1 0 36966 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_78_385
timestamp 1607639953
transform 1 0 36506 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1607639953
transform 1 0 36690 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_410
timestamp 1607639953
transform 1 0 38806 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_398
timestamp 1607639953
transform 1 0 37702 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1000
timestamp 1607639953
transform 1 0 37610 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_434
timestamp 1607639953
transform 1 0 41014 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_422
timestamp 1607639953
transform 1 0 39910 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_459
timestamp 1607639953
transform 1 0 43314 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_446
timestamp 1607639953
transform 1 0 42118 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1001
timestamp 1607639953
transform 1 0 43222 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_483
timestamp 1607639953
transform 1 0 45522 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_471
timestamp 1607639953
transform 1 0 44418 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_495
timestamp 1607639953
transform 1 0 46626 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_520
timestamp 1607639953
transform 1 0 48926 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_507
timestamp 1607639953
transform 1 0 47730 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1002
timestamp 1607639953
transform 1 0 48834 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_544
timestamp 1607639953
transform 1 0 51134 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_532
timestamp 1607639953
transform 1 0 50030 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_568
timestamp 1607639953
transform 1 0 53342 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_556
timestamp 1607639953
transform 1 0 52238 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_593
timestamp 1607639953
transform 1 0 55642 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_581
timestamp 1607639953
transform 1 0 54538 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1003
timestamp 1607639953
transform 1 0 54446 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_605
timestamp 1607639953
transform 1 0 56746 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_617
timestamp 1607639953
transform 1 0 57850 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1607639953
transform -1 0 58862 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_20
timestamp 1607639953
transform 1 0 2926 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_15
timestamp 1607639953
transform 1 0 2466 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1607639953
transform 1 0 1362 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1607639953
transform 1 0 2466 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1607639953
transform 1 0 1362 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1607639953
transform 1 0 1086 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1607639953
transform 1 0 1086 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _077_
timestamp 1607639953
transform 1 0 2650 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_44
timestamp 1607639953
transform 1 0 5134 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_32
timestamp 1607639953
transform 1 0 4030 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_28
timestamp 1607639953
transform 1 0 3662 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1607639953
transform 1 0 4674 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1607639953
transform 1 0 3570 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1014
timestamp 1607639953
transform 1 0 3938 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_56
timestamp 1607639953
transform 1 0 6238 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_62
timestamp 1607639953
transform 1 0 6790 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_59
timestamp 1607639953
transform 1 0 6514 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_51
timestamp 1607639953
transform 1 0 5778 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1004
timestamp 1607639953
transform 1 0 6698 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_80
timestamp 1607639953
transform 1 0 8446 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_68
timestamp 1607639953
transform 1 0 7342 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_86
timestamp 1607639953
transform 1 0 8998 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_74
timestamp 1607639953
transform 1 0 7894 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _124_
timestamp 1607639953
transform 1 0 8998 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_105
timestamp 1607639953
transform 1 0 10746 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_93
timestamp 1607639953
transform 1 0 9642 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_89
timestamp 1607639953
transform 1 0 9274 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_110
timestamp 1607639953
transform 1 0 11206 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_98
timestamp 1607639953
transform 1 0 10102 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1015
timestamp 1607639953
transform 1 0 9550 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_129
timestamp 1607639953
transform 1 0 12954 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_117
timestamp 1607639953
transform 1 0 11850 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_123
timestamp 1607639953
transform 1 0 12402 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1005
timestamp 1607639953
transform 1 0 12310 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_154
timestamp 1607639953
transform 1 0 15254 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_141
timestamp 1607639953
transform 1 0 14058 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_147
timestamp 1607639953
transform 1 0 14610 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_135
timestamp 1607639953
transform 1 0 13506 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1016
timestamp 1607639953
transform 1 0 15162 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_166
timestamp 1607639953
transform 1 0 16358 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_171
timestamp 1607639953
transform 1 0 16818 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_159
timestamp 1607639953
transform 1 0 15714 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_190
timestamp 1607639953
transform 1 0 18566 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_178
timestamp 1607639953
transform 1 0 17462 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_196
timestamp 1607639953
transform 1 0 19118 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_184
timestamp 1607639953
transform 1 0 18014 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1006
timestamp 1607639953
transform 1 0 17922 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_215
timestamp 1607639953
transform 1 0 20866 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_212
timestamp 1607639953
transform 1 0 20590 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_208
timestamp 1607639953
transform 1 0 20222 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_202
timestamp 1607639953
transform 1 0 19670 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_217
timestamp 1607639953
transform 1 0 21050 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_208
timestamp 1607639953
transform 1 0 20222 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1017
timestamp 1607639953
transform 1 0 20774 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _196_
timestamp 1607639953
transform 1 0 20774 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _191_
timestamp 1607639953
transform 1 0 20314 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_239
timestamp 1607639953
transform 1 0 23074 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_227
timestamp 1607639953
transform 1 0 21970 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_241
timestamp 1607639953
transform 1 0 23258 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_229
timestamp 1607639953
transform 1 0 22154 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_263
timestamp 1607639953
transform 1 0 25282 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_251
timestamp 1607639953
transform 1 0 24178 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_257
timestamp 1607639953
transform 1 0 24730 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_245
timestamp 1607639953
transform 1 0 23626 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1007
timestamp 1607639953
transform 1 0 23534 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_276
timestamp 1607639953
transform 1 0 26478 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1607639953
transform 1 0 26938 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_269
timestamp 1607639953
transform 1 0 25834 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1018
timestamp 1607639953
transform 1 0 26386 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_300
timestamp 1607639953
transform 1 0 28686 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_288
timestamp 1607639953
transform 1 0 27582 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1607639953
transform 1 0 28042 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1008
timestamp 1607639953
transform 1 0 29146 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _117_
timestamp 1607639953
transform 1 0 29238 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_324
timestamp 1607639953
transform 1 0 30894 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_312
timestamp 1607639953
transform 1 0 29790 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_321
timestamp 1607639953
transform 1 0 30618 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_309
timestamp 1607639953
transform 1 0 29514 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_347
timestamp 1607639953
transform 1 0 33010 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_343
timestamp 1607639953
transform 1 0 32642 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_337
timestamp 1607639953
transform 1 0 32090 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_345
timestamp 1607639953
transform 1 0 32826 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_333
timestamp 1607639953
transform 1 0 31722 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1019
timestamp 1607639953
transform 1 0 31998 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _078_
timestamp 1607639953
transform 1 0 32734 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_371
timestamp 1607639953
transform 1 0 35218 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_359
timestamp 1607639953
transform 1 0 34114 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_367
timestamp 1607639953
transform 1 0 34850 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_365
timestamp 1607639953
transform 1 0 34666 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_357
timestamp 1607639953
transform 1 0 33930 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1009
timestamp 1607639953
transform 1 0 34758 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_395
timestamp 1607639953
transform 1 0 37426 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_383
timestamp 1607639953
transform 1 0 36322 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_391
timestamp 1607639953
transform 1 0 37058 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_379
timestamp 1607639953
transform 1 0 35954 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_410
timestamp 1607639953
transform 1 0 38806 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_398
timestamp 1607639953
transform 1 0 37702 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_413
timestamp 1607639953
transform 1 0 39082 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_409
timestamp 1607639953
transform 1 0 38714 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_403
timestamp 1607639953
transform 1 0 38162 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1020
timestamp 1607639953
transform 1 0 37610 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1607639953
transform 1 0 38806 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_434
timestamp 1607639953
transform 1 0 41014 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_422
timestamp 1607639953
transform 1 0 39910 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_440
timestamp 1607639953
transform 1 0 41566 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_428
timestamp 1607639953
transform 1 0 40462 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_425
timestamp 1607639953
transform 1 0 40186 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1010
timestamp 1607639953
transform 1 0 40370 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_459
timestamp 1607639953
transform 1 0 43314 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_446
timestamp 1607639953
transform 1 0 42118 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_452
timestamp 1607639953
transform 1 0 42670 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1021
timestamp 1607639953
transform 1 0 43222 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_483
timestamp 1607639953
transform 1 0 45522 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_471
timestamp 1607639953
transform 1 0 44418 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_476
timestamp 1607639953
transform 1 0 44878 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_464
timestamp 1607639953
transform 1 0 43774 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_495
timestamp 1607639953
transform 1 0 46626 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_501
timestamp 1607639953
transform 1 0 47178 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_489
timestamp 1607639953
transform 1 0 46074 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1011
timestamp 1607639953
transform 1 0 45982 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_520
timestamp 1607639953
transform 1 0 48926 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_507
timestamp 1607639953
transform 1 0 47730 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_525
timestamp 1607639953
transform 1 0 49386 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_513
timestamp 1607639953
transform 1 0 48282 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1022
timestamp 1607639953
transform 1 0 48834 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_544
timestamp 1607639953
transform 1 0 51134 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_532
timestamp 1607639953
transform 1 0 50030 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_550
timestamp 1607639953
transform 1 0 51686 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_537
timestamp 1607639953
transform 1 0 50490 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1012
timestamp 1607639953
transform 1 0 51594 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_568
timestamp 1607639953
transform 1 0 53342 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_556
timestamp 1607639953
transform 1 0 52238 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_562
timestamp 1607639953
transform 1 0 52790 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_593
timestamp 1607639953
transform 1 0 55642 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_581
timestamp 1607639953
transform 1 0 54538 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_586
timestamp 1607639953
transform 1 0 54998 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_574
timestamp 1607639953
transform 1 0 53894 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1023
timestamp 1607639953
transform 1 0 54446 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_605
timestamp 1607639953
transform 1 0 56746 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_611
timestamp 1607639953
transform 1 0 57298 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_598
timestamp 1607639953
transform 1 0 56102 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1013
timestamp 1607639953
transform 1 0 57206 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_617
timestamp 1607639953
transform 1 0 57850 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_623
timestamp 1607639953
transform 1 0 58402 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1607639953
transform -1 0 58862 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1607639953
transform -1 0 58862 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1607639953
transform 1 0 2466 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1607639953
transform 1 0 1362 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1607639953
transform 1 0 1086 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_39
timestamp 1607639953
transform 1 0 4674 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1607639953
transform 1 0 3570 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_62
timestamp 1607639953
transform 1 0 6790 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_59
timestamp 1607639953
transform 1 0 6514 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_51
timestamp 1607639953
transform 1 0 5778 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1024
timestamp 1607639953
transform 1 0 6698 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_86
timestamp 1607639953
transform 1 0 8998 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_74
timestamp 1607639953
transform 1 0 7894 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_110
timestamp 1607639953
transform 1 0 11206 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_98
timestamp 1607639953
transform 1 0 10102 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_123
timestamp 1607639953
transform 1 0 12402 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1025
timestamp 1607639953
transform 1 0 12310 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_147
timestamp 1607639953
transform 1 0 14610 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_135
timestamp 1607639953
transform 1 0 13506 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_171
timestamp 1607639953
transform 1 0 16818 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_159
timestamp 1607639953
transform 1 0 15714 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_196
timestamp 1607639953
transform 1 0 19118 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_184
timestamp 1607639953
transform 1 0 18014 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1026
timestamp 1607639953
transform 1 0 17922 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_220
timestamp 1607639953
transform 1 0 21326 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_208
timestamp 1607639953
transform 1 0 20222 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_232
timestamp 1607639953
transform 1 0 22430 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_257
timestamp 1607639953
transform 1 0 24730 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_245
timestamp 1607639953
transform 1 0 23626 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1027
timestamp 1607639953
transform 1 0 23534 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1607639953
transform 1 0 26938 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_269
timestamp 1607639953
transform 1 0 25834 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_306
timestamp 1607639953
transform 1 0 29238 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1607639953
transform 1 0 28042 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1028
timestamp 1607639953
transform 1 0 29146 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_330
timestamp 1607639953
transform 1 0 31446 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_318
timestamp 1607639953
transform 1 0 30342 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_350
timestamp 1607639953
transform 1 0 33286 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_342
timestamp 1607639953
transform 1 0 32550 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_367
timestamp 1607639953
transform 1 0 34850 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_364
timestamp 1607639953
transform 1 0 34574 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_356
timestamp 1607639953
transform 1 0 33838 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1029
timestamp 1607639953
transform 1 0 34758 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1607639953
transform 1 0 33562 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_391
timestamp 1607639953
transform 1 0 37058 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_379
timestamp 1607639953
transform 1 0 35954 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_415
timestamp 1607639953
transform 1 0 39266 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_403
timestamp 1607639953
transform 1 0 38162 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_440
timestamp 1607639953
transform 1 0 41566 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_428
timestamp 1607639953
transform 1 0 40462 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1030
timestamp 1607639953
transform 1 0 40370 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_452
timestamp 1607639953
transform 1 0 42670 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_476
timestamp 1607639953
transform 1 0 44878 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_464
timestamp 1607639953
transform 1 0 43774 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_501
timestamp 1607639953
transform 1 0 47178 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_489
timestamp 1607639953
transform 1 0 46074 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1031
timestamp 1607639953
transform 1 0 45982 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_525
timestamp 1607639953
transform 1 0 49386 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_513
timestamp 1607639953
transform 1 0 48282 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_509
timestamp 1607639953
transform 1 0 47914 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _016_
timestamp 1607639953
transform 1 0 48006 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_550
timestamp 1607639953
transform 1 0 51686 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_537
timestamp 1607639953
transform 1 0 50490 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1032
timestamp 1607639953
transform 1 0 51594 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_562
timestamp 1607639953
transform 1 0 52790 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_586
timestamp 1607639953
transform 1 0 54998 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_574
timestamp 1607639953
transform 1 0 53894 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_611
timestamp 1607639953
transform 1 0 57298 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_598
timestamp 1607639953
transform 1 0 56102 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1033
timestamp 1607639953
transform 1 0 57206 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_624
timestamp 1607639953
transform 1 0 58494 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_619
timestamp 1607639953
transform 1 0 58034 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1607639953
transform -1 0 58862 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _158_
timestamp 1607639953
transform 1 0 58218 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1607639953
transform 1 0 2466 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1607639953
transform 1 0 1362 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1607639953
transform 1 0 1086 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_44
timestamp 1607639953
transform 1 0 5134 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_32
timestamp 1607639953
transform 1 0 4030 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_27
timestamp 1607639953
transform 1 0 3570 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1034
timestamp 1607639953
transform 1 0 3938 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_56
timestamp 1607639953
transform 1 0 6238 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_80
timestamp 1607639953
transform 1 0 8446 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_68
timestamp 1607639953
transform 1 0 7342 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_105
timestamp 1607639953
transform 1 0 10746 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_93
timestamp 1607639953
transform 1 0 9642 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1035
timestamp 1607639953
transform 1 0 9550 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_129
timestamp 1607639953
transform 1 0 12954 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_117
timestamp 1607639953
transform 1 0 11850 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_154
timestamp 1607639953
transform 1 0 15254 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_141
timestamp 1607639953
transform 1 0 14058 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1036
timestamp 1607639953
transform 1 0 15162 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_166
timestamp 1607639953
transform 1 0 16358 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_190
timestamp 1607639953
transform 1 0 18566 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_178
timestamp 1607639953
transform 1 0 17462 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_215
timestamp 1607639953
transform 1 0 20866 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_202
timestamp 1607639953
transform 1 0 19670 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1037
timestamp 1607639953
transform 1 0 20774 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_239
timestamp 1607639953
transform 1 0 23074 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_227
timestamp 1607639953
transform 1 0 21970 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_263
timestamp 1607639953
transform 1 0 25282 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_251
timestamp 1607639953
transform 1 0 24178 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_276
timestamp 1607639953
transform 1 0 26478 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1038
timestamp 1607639953
transform 1 0 26386 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_300
timestamp 1607639953
transform 1 0 28686 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_288
timestamp 1607639953
transform 1 0 27582 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_324
timestamp 1607639953
transform 1 0 30894 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_312
timestamp 1607639953
transform 1 0 29790 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_349
timestamp 1607639953
transform 1 0 33194 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1607639953
transform 1 0 32090 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1039
timestamp 1607639953
transform 1 0 31998 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_371
timestamp 1607639953
transform 1 0 35218 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_359
timestamp 1607639953
transform 1 0 34114 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_355
timestamp 1607639953
transform 1 0 33746 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1607639953
transform 1 0 33838 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_395
timestamp 1607639953
transform 1 0 37426 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_383
timestamp 1607639953
transform 1 0 36322 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_410
timestamp 1607639953
transform 1 0 38806 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_398
timestamp 1607639953
transform 1 0 37702 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1040
timestamp 1607639953
transform 1 0 37610 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_434
timestamp 1607639953
transform 1 0 41014 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_422
timestamp 1607639953
transform 1 0 39910 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_459
timestamp 1607639953
transform 1 0 43314 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_446
timestamp 1607639953
transform 1 0 42118 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1041
timestamp 1607639953
transform 1 0 43222 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_483
timestamp 1607639953
transform 1 0 45522 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_471
timestamp 1607639953
transform 1 0 44418 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_495
timestamp 1607639953
transform 1 0 46626 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_520
timestamp 1607639953
transform 1 0 48926 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_507
timestamp 1607639953
transform 1 0 47730 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1042
timestamp 1607639953
transform 1 0 48834 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_544
timestamp 1607639953
transform 1 0 51134 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_532
timestamp 1607639953
transform 1 0 50030 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_568
timestamp 1607639953
transform 1 0 53342 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_556
timestamp 1607639953
transform 1 0 52238 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_593
timestamp 1607639953
transform 1 0 55642 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_581
timestamp 1607639953
transform 1 0 54538 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1043
timestamp 1607639953
transform 1 0 54446 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_605
timestamp 1607639953
transform 1 0 56746 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_617
timestamp 1607639953
transform 1 0 57850 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1607639953
transform -1 0 58862 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_15
timestamp 1607639953
transform 1 0 2466 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_3
timestamp 1607639953
transform 1 0 1362 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1607639953
transform 1 0 1086 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_39
timestamp 1607639953
transform 1 0 4674 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_27
timestamp 1607639953
transform 1 0 3570 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_62
timestamp 1607639953
transform 1 0 6790 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_59
timestamp 1607639953
transform 1 0 6514 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_83_51
timestamp 1607639953
transform 1 0 5778 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1044
timestamp 1607639953
transform 1 0 6698 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_86
timestamp 1607639953
transform 1 0 8998 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_74
timestamp 1607639953
transform 1 0 7894 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_110
timestamp 1607639953
transform 1 0 11206 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_98
timestamp 1607639953
transform 1 0 10102 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_123
timestamp 1607639953
transform 1 0 12402 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1045
timestamp 1607639953
transform 1 0 12310 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_147
timestamp 1607639953
transform 1 0 14610 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_135
timestamp 1607639953
transform 1 0 13506 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_171
timestamp 1607639953
transform 1 0 16818 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_159
timestamp 1607639953
transform 1 0 15714 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_196
timestamp 1607639953
transform 1 0 19118 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_184
timestamp 1607639953
transform 1 0 18014 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1046
timestamp 1607639953
transform 1 0 17922 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_220
timestamp 1607639953
transform 1 0 21326 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_208
timestamp 1607639953
transform 1 0 20222 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_232
timestamp 1607639953
transform 1 0 22430 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_257
timestamp 1607639953
transform 1 0 24730 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_245
timestamp 1607639953
transform 1 0 23626 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1047
timestamp 1607639953
transform 1 0 23534 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_281
timestamp 1607639953
transform 1 0 26938 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_269
timestamp 1607639953
transform 1 0 25834 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_306
timestamp 1607639953
transform 1 0 29238 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_293
timestamp 1607639953
transform 1 0 28042 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1048
timestamp 1607639953
transform 1 0 29146 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_330
timestamp 1607639953
transform 1 0 31446 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_318
timestamp 1607639953
transform 1 0 30342 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_342
timestamp 1607639953
transform 1 0 32550 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_367
timestamp 1607639953
transform 1 0 34850 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_354
timestamp 1607639953
transform 1 0 33654 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1049
timestamp 1607639953
transform 1 0 34758 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_391
timestamp 1607639953
transform 1 0 37058 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_379
timestamp 1607639953
transform 1 0 35954 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_415
timestamp 1607639953
transform 1 0 39266 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_403
timestamp 1607639953
transform 1 0 38162 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_440
timestamp 1607639953
transform 1 0 41566 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_428
timestamp 1607639953
transform 1 0 40462 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1050
timestamp 1607639953
transform 1 0 40370 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_452
timestamp 1607639953
transform 1 0 42670 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_476
timestamp 1607639953
transform 1 0 44878 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_464
timestamp 1607639953
transform 1 0 43774 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_501
timestamp 1607639953
transform 1 0 47178 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_489
timestamp 1607639953
transform 1 0 46074 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1051
timestamp 1607639953
transform 1 0 45982 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_525
timestamp 1607639953
transform 1 0 49386 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_513
timestamp 1607639953
transform 1 0 48282 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_550
timestamp 1607639953
transform 1 0 51686 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_537
timestamp 1607639953
transform 1 0 50490 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1052
timestamp 1607639953
transform 1 0 51594 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_562
timestamp 1607639953
transform 1 0 52790 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_586
timestamp 1607639953
transform 1 0 54998 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_574
timestamp 1607639953
transform 1 0 53894 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_611
timestamp 1607639953
transform 1 0 57298 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_598
timestamp 1607639953
transform 1 0 56102 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1053
timestamp 1607639953
transform 1 0 57206 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_623
timestamp 1607639953
transform 1 0 58402 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1607639953
transform -1 0 58862 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_15
timestamp 1607639953
transform 1 0 2466 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_3
timestamp 1607639953
transform 1 0 1362 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1607639953
transform 1 0 1086 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_44
timestamp 1607639953
transform 1 0 5134 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_32
timestamp 1607639953
transform 1 0 4030 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_27
timestamp 1607639953
transform 1 0 3570 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1054
timestamp 1607639953
transform 1 0 3938 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_56
timestamp 1607639953
transform 1 0 6238 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_80
timestamp 1607639953
transform 1 0 8446 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_68
timestamp 1607639953
transform 1 0 7342 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_105
timestamp 1607639953
transform 1 0 10746 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_93
timestamp 1607639953
transform 1 0 9642 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1055
timestamp 1607639953
transform 1 0 9550 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_129
timestamp 1607639953
transform 1 0 12954 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_117
timestamp 1607639953
transform 1 0 11850 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_154
timestamp 1607639953
transform 1 0 15254 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_141
timestamp 1607639953
transform 1 0 14058 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1056
timestamp 1607639953
transform 1 0 15162 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_166
timestamp 1607639953
transform 1 0 16358 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_190
timestamp 1607639953
transform 1 0 18566 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_178
timestamp 1607639953
transform 1 0 17462 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_215
timestamp 1607639953
transform 1 0 20866 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_202
timestamp 1607639953
transform 1 0 19670 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1057
timestamp 1607639953
transform 1 0 20774 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_239
timestamp 1607639953
transform 1 0 23074 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_227
timestamp 1607639953
transform 1 0 21970 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_263
timestamp 1607639953
transform 1 0 25282 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_251
timestamp 1607639953
transform 1 0 24178 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_276
timestamp 1607639953
transform 1 0 26478 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1058
timestamp 1607639953
transform 1 0 26386 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_300
timestamp 1607639953
transform 1 0 28686 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_288
timestamp 1607639953
transform 1 0 27582 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_324
timestamp 1607639953
transform 1 0 30894 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_312
timestamp 1607639953
transform 1 0 29790 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_349
timestamp 1607639953
transform 1 0 33194 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_337
timestamp 1607639953
transform 1 0 32090 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1059
timestamp 1607639953
transform 1 0 31998 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_373
timestamp 1607639953
transform 1 0 35402 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_361
timestamp 1607639953
transform 1 0 34298 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_385
timestamp 1607639953
transform 1 0 36506 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_410
timestamp 1607639953
transform 1 0 38806 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_398
timestamp 1607639953
transform 1 0 37702 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1060
timestamp 1607639953
transform 1 0 37610 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_434
timestamp 1607639953
transform 1 0 41014 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_422
timestamp 1607639953
transform 1 0 39910 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_459
timestamp 1607639953
transform 1 0 43314 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_446
timestamp 1607639953
transform 1 0 42118 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1061
timestamp 1607639953
transform 1 0 43222 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_483
timestamp 1607639953
transform 1 0 45522 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_471
timestamp 1607639953
transform 1 0 44418 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_497
timestamp 1607639953
transform 1 0 46810 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_491
timestamp 1607639953
transform 1 0 46258 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _102_
timestamp 1607639953
transform 1 0 46534 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_520
timestamp 1607639953
transform 1 0 48926 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_84_517
timestamp 1607639953
transform 1 0 48650 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_84_509
timestamp 1607639953
transform 1 0 47914 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1062
timestamp 1607639953
transform 1 0 48834 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_544
timestamp 1607639953
transform 1 0 51134 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_532
timestamp 1607639953
transform 1 0 50030 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_568
timestamp 1607639953
transform 1 0 53342 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_556
timestamp 1607639953
transform 1 0 52238 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_593
timestamp 1607639953
transform 1 0 55642 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_581
timestamp 1607639953
transform 1 0 54538 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1063
timestamp 1607639953
transform 1 0 54446 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_605
timestamp 1607639953
transform 1 0 56746 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_617
timestamp 1607639953
transform 1 0 57850 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1607639953
transform -1 0 58862 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_15
timestamp 1607639953
transform 1 0 2466 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_3
timestamp 1607639953
transform 1 0 1362 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1607639953
transform 1 0 2466 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1607639953
transform 1 0 1362 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1607639953
transform 1 0 1086 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1607639953
transform 1 0 1086 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_44
timestamp 1607639953
transform 1 0 5134 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_32
timestamp 1607639953
transform 1 0 4030 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_27
timestamp 1607639953
transform 1 0 3570 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_39
timestamp 1607639953
transform 1 0 4674 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1607639953
transform 1 0 3570 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1074
timestamp 1607639953
transform 1 0 3938 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_56
timestamp 1607639953
transform 1 0 6238 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_62
timestamp 1607639953
transform 1 0 6790 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_59
timestamp 1607639953
transform 1 0 6514 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_85_51
timestamp 1607639953
transform 1 0 5778 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1064
timestamp 1607639953
transform 1 0 6698 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_80
timestamp 1607639953
transform 1 0 8446 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_68
timestamp 1607639953
transform 1 0 7342 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_86
timestamp 1607639953
transform 1 0 8998 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_74
timestamp 1607639953
transform 1 0 7894 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_105
timestamp 1607639953
transform 1 0 10746 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_93
timestamp 1607639953
transform 1 0 9642 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_110
timestamp 1607639953
transform 1 0 11206 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_98
timestamp 1607639953
transform 1 0 10102 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1075
timestamp 1607639953
transform 1 0 9550 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_129
timestamp 1607639953
transform 1 0 12954 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_117
timestamp 1607639953
transform 1 0 11850 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_123
timestamp 1607639953
transform 1 0 12402 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1065
timestamp 1607639953
transform 1 0 12310 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_154
timestamp 1607639953
transform 1 0 15254 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_141
timestamp 1607639953
transform 1 0 14058 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_147
timestamp 1607639953
transform 1 0 14610 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_135
timestamp 1607639953
transform 1 0 13506 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1076
timestamp 1607639953
transform 1 0 15162 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_166
timestamp 1607639953
transform 1 0 16358 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_171
timestamp 1607639953
transform 1 0 16818 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_159
timestamp 1607639953
transform 1 0 15714 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_190
timestamp 1607639953
transform 1 0 18566 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_178
timestamp 1607639953
transform 1 0 17462 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_196
timestamp 1607639953
transform 1 0 19118 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_184
timestamp 1607639953
transform 1 0 18014 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1066
timestamp 1607639953
transform 1 0 17922 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_215
timestamp 1607639953
transform 1 0 20866 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_202
timestamp 1607639953
transform 1 0 19670 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_220
timestamp 1607639953
transform 1 0 21326 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_208
timestamp 1607639953
transform 1 0 20222 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1077
timestamp 1607639953
transform 1 0 20774 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_239
timestamp 1607639953
transform 1 0 23074 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_227
timestamp 1607639953
transform 1 0 21970 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_240
timestamp 1607639953
transform 1 0 23166 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_236
timestamp 1607639953
transform 1 0 22798 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_232
timestamp 1607639953
transform 1 0 22430 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1607639953
transform 1 0 22890 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_263
timestamp 1607639953
transform 1 0 25282 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_251
timestamp 1607639953
transform 1 0 24178 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_257
timestamp 1607639953
transform 1 0 24730 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_245
timestamp 1607639953
transform 1 0 23626 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1067
timestamp 1607639953
transform 1 0 23534 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_276
timestamp 1607639953
transform 1 0 26478 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_281
timestamp 1607639953
transform 1 0 26938 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_269
timestamp 1607639953
transform 1 0 25834 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1078
timestamp 1607639953
transform 1 0 26386 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_300
timestamp 1607639953
transform 1 0 28686 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_288
timestamp 1607639953
transform 1 0 27582 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_306
timestamp 1607639953
transform 1 0 29238 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_293
timestamp 1607639953
transform 1 0 28042 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1068
timestamp 1607639953
transform 1 0 29146 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_324
timestamp 1607639953
transform 1 0 30894 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_312
timestamp 1607639953
transform 1 0 29790 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_330
timestamp 1607639953
transform 1 0 31446 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_318
timestamp 1607639953
transform 1 0 30342 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_349
timestamp 1607639953
transform 1 0 33194 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_337
timestamp 1607639953
transform 1 0 32090 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_342
timestamp 1607639953
transform 1 0 32550 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1079
timestamp 1607639953
transform 1 0 31998 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_373
timestamp 1607639953
transform 1 0 35402 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_361
timestamp 1607639953
transform 1 0 34298 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_367
timestamp 1607639953
transform 1 0 34850 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_365
timestamp 1607639953
transform 1 0 34666 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_85_359
timestamp 1607639953
transform 1 0 34114 0 1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_85_354
timestamp 1607639953
transform 1 0 33654 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1069
timestamp 1607639953
transform 1 0 34758 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _131_
timestamp 1607639953
transform 1 0 33838 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_385
timestamp 1607639953
transform 1 0 36506 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_391
timestamp 1607639953
transform 1 0 37058 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_379
timestamp 1607639953
transform 1 0 35954 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_410
timestamp 1607639953
transform 1 0 38806 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_398
timestamp 1607639953
transform 1 0 37702 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_415
timestamp 1607639953
transform 1 0 39266 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_403
timestamp 1607639953
transform 1 0 38162 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1080
timestamp 1607639953
transform 1 0 37610 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_434
timestamp 1607639953
transform 1 0 41014 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_422
timestamp 1607639953
transform 1 0 39910 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_440
timestamp 1607639953
transform 1 0 41566 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_428
timestamp 1607639953
transform 1 0 40462 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1070
timestamp 1607639953
transform 1 0 40370 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_459
timestamp 1607639953
transform 1 0 43314 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_446
timestamp 1607639953
transform 1 0 42118 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_452
timestamp 1607639953
transform 1 0 42670 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1081
timestamp 1607639953
transform 1 0 43222 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_483
timestamp 1607639953
transform 1 0 45522 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_471
timestamp 1607639953
transform 1 0 44418 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_476
timestamp 1607639953
transform 1 0 44878 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_464
timestamp 1607639953
transform 1 0 43774 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_495
timestamp 1607639953
transform 1 0 46626 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_501
timestamp 1607639953
transform 1 0 47178 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_489
timestamp 1607639953
transform 1 0 46074 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1071
timestamp 1607639953
transform 1 0 45982 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_520
timestamp 1607639953
transform 1 0 48926 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_518
timestamp 1607639953
transform 1 0 48742 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_507
timestamp 1607639953
transform 1 0 47730 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_525
timestamp 1607639953
transform 1 0 49386 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_513
timestamp 1607639953
transform 1 0 48282 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1082
timestamp 1607639953
transform 1 0 48834 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _070_
timestamp 1607639953
transform 1 0 48466 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_544
timestamp 1607639953
transform 1 0 51134 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_532
timestamp 1607639953
transform 1 0 50030 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_550
timestamp 1607639953
transform 1 0 51686 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_537
timestamp 1607639953
transform 1 0 50490 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1072
timestamp 1607639953
transform 1 0 51594 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_568
timestamp 1607639953
transform 1 0 53342 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_556
timestamp 1607639953
transform 1 0 52238 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_562
timestamp 1607639953
transform 1 0 52790 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_593
timestamp 1607639953
transform 1 0 55642 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_581
timestamp 1607639953
transform 1 0 54538 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_586
timestamp 1607639953
transform 1 0 54998 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_574
timestamp 1607639953
transform 1 0 53894 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1083
timestamp 1607639953
transform 1 0 54446 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_605
timestamp 1607639953
transform 1 0 56746 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_611
timestamp 1607639953
transform 1 0 57298 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_598
timestamp 1607639953
transform 1 0 56102 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1073
timestamp 1607639953
transform 1 0 57206 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_617
timestamp 1607639953
transform 1 0 57850 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_623
timestamp 1607639953
transform 1 0 58402 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1607639953
transform -1 0 58862 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1607639953
transform -1 0 58862 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_15
timestamp 1607639953
transform 1 0 2466 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_3
timestamp 1607639953
transform 1 0 1362 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1607639953
transform 1 0 1086 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_39
timestamp 1607639953
transform 1 0 4674 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_27
timestamp 1607639953
transform 1 0 3570 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_62
timestamp 1607639953
transform 1 0 6790 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_59
timestamp 1607639953
transform 1 0 6514 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_87_51
timestamp 1607639953
transform 1 0 5778 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1084
timestamp 1607639953
transform 1 0 6698 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_86
timestamp 1607639953
transform 1 0 8998 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_74
timestamp 1607639953
transform 1 0 7894 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_110
timestamp 1607639953
transform 1 0 11206 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_98
timestamp 1607639953
transform 1 0 10102 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_123
timestamp 1607639953
transform 1 0 12402 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1085
timestamp 1607639953
transform 1 0 12310 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_147
timestamp 1607639953
transform 1 0 14610 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_135
timestamp 1607639953
transform 1 0 13506 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_171
timestamp 1607639953
transform 1 0 16818 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_159
timestamp 1607639953
transform 1 0 15714 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_196
timestamp 1607639953
transform 1 0 19118 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_184
timestamp 1607639953
transform 1 0 18014 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1086
timestamp 1607639953
transform 1 0 17922 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_220
timestamp 1607639953
transform 1 0 21326 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_208
timestamp 1607639953
transform 1 0 20222 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_232
timestamp 1607639953
transform 1 0 22430 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_257
timestamp 1607639953
transform 1 0 24730 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_245
timestamp 1607639953
transform 1 0 23626 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1087
timestamp 1607639953
transform 1 0 23534 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_281
timestamp 1607639953
transform 1 0 26938 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_269
timestamp 1607639953
transform 1 0 25834 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_306
timestamp 1607639953
transform 1 0 29238 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_293
timestamp 1607639953
transform 1 0 28042 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1088
timestamp 1607639953
transform 1 0 29146 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_330
timestamp 1607639953
transform 1 0 31446 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_318
timestamp 1607639953
transform 1 0 30342 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_342
timestamp 1607639953
transform 1 0 32550 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_367
timestamp 1607639953
transform 1 0 34850 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_87_365
timestamp 1607639953
transform 1 0 34666 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_357
timestamp 1607639953
transform 1 0 33930 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1089
timestamp 1607639953
transform 1 0 34758 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1607639953
transform 1 0 33654 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_391
timestamp 1607639953
transform 1 0 37058 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_379
timestamp 1607639953
transform 1 0 35954 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_415
timestamp 1607639953
transform 1 0 39266 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_403
timestamp 1607639953
transform 1 0 38162 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_440
timestamp 1607639953
transform 1 0 41566 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_428
timestamp 1607639953
transform 1 0 40462 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1090
timestamp 1607639953
transform 1 0 40370 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_452
timestamp 1607639953
transform 1 0 42670 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_476
timestamp 1607639953
transform 1 0 44878 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_464
timestamp 1607639953
transform 1 0 43774 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_501
timestamp 1607639953
transform 1 0 47178 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_489
timestamp 1607639953
transform 1 0 46074 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1091
timestamp 1607639953
transform 1 0 45982 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_525
timestamp 1607639953
transform 1 0 49386 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_513
timestamp 1607639953
transform 1 0 48282 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_550
timestamp 1607639953
transform 1 0 51686 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_537
timestamp 1607639953
transform 1 0 50490 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1092
timestamp 1607639953
transform 1 0 51594 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_562
timestamp 1607639953
transform 1 0 52790 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_586
timestamp 1607639953
transform 1 0 54998 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_574
timestamp 1607639953
transform 1 0 53894 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_611
timestamp 1607639953
transform 1 0 57298 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_598
timestamp 1607639953
transform 1 0 56102 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1093
timestamp 1607639953
transform 1 0 57206 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_623
timestamp 1607639953
transform 1 0 58402 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1607639953
transform -1 0 58862 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_15
timestamp 1607639953
transform 1 0 2466 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_3
timestamp 1607639953
transform 1 0 1362 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1607639953
transform 1 0 1086 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_44
timestamp 1607639953
transform 1 0 5134 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_32
timestamp 1607639953
transform 1 0 4030 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_27
timestamp 1607639953
transform 1 0 3570 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1094
timestamp 1607639953
transform 1 0 3938 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_56
timestamp 1607639953
transform 1 0 6238 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_80
timestamp 1607639953
transform 1 0 8446 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_68
timestamp 1607639953
transform 1 0 7342 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_105
timestamp 1607639953
transform 1 0 10746 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_93
timestamp 1607639953
transform 1 0 9642 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1095
timestamp 1607639953
transform 1 0 9550 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_129
timestamp 1607639953
transform 1 0 12954 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_117
timestamp 1607639953
transform 1 0 11850 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_154
timestamp 1607639953
transform 1 0 15254 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_141
timestamp 1607639953
transform 1 0 14058 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1096
timestamp 1607639953
transform 1 0 15162 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_166
timestamp 1607639953
transform 1 0 16358 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_190
timestamp 1607639953
transform 1 0 18566 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_178
timestamp 1607639953
transform 1 0 17462 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_215
timestamp 1607639953
transform 1 0 20866 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_202
timestamp 1607639953
transform 1 0 19670 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1097
timestamp 1607639953
transform 1 0 20774 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_239
timestamp 1607639953
transform 1 0 23074 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_227
timestamp 1607639953
transform 1 0 21970 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_263
timestamp 1607639953
transform 1 0 25282 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_251
timestamp 1607639953
transform 1 0 24178 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_276
timestamp 1607639953
transform 1 0 26478 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1098
timestamp 1607639953
transform 1 0 26386 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_300
timestamp 1607639953
transform 1 0 28686 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_288
timestamp 1607639953
transform 1 0 27582 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_324
timestamp 1607639953
transform 1 0 30894 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_312
timestamp 1607639953
transform 1 0 29790 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_349
timestamp 1607639953
transform 1 0 33194 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_337
timestamp 1607639953
transform 1 0 32090 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1099
timestamp 1607639953
transform 1 0 31998 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_373
timestamp 1607639953
transform 1 0 35402 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_361
timestamp 1607639953
transform 1 0 34298 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_385
timestamp 1607639953
transform 1 0 36506 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_410
timestamp 1607639953
transform 1 0 38806 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_398
timestamp 1607639953
transform 1 0 37702 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1100
timestamp 1607639953
transform 1 0 37610 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_434
timestamp 1607639953
transform 1 0 41014 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_422
timestamp 1607639953
transform 1 0 39910 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_459
timestamp 1607639953
transform 1 0 43314 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_446
timestamp 1607639953
transform 1 0 42118 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1101
timestamp 1607639953
transform 1 0 43222 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_483
timestamp 1607639953
transform 1 0 45522 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_471
timestamp 1607639953
transform 1 0 44418 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_495
timestamp 1607639953
transform 1 0 46626 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_520
timestamp 1607639953
transform 1 0 48926 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_507
timestamp 1607639953
transform 1 0 47730 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1102
timestamp 1607639953
transform 1 0 48834 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_544
timestamp 1607639953
transform 1 0 51134 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_532
timestamp 1607639953
transform 1 0 50030 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_568
timestamp 1607639953
transform 1 0 53342 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_556
timestamp 1607639953
transform 1 0 52238 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_593
timestamp 1607639953
transform 1 0 55642 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_581
timestamp 1607639953
transform 1 0 54538 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1103
timestamp 1607639953
transform 1 0 54446 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_605
timestamp 1607639953
transform 1 0 56746 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_617
timestamp 1607639953
transform 1 0 57850 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1607639953
transform -1 0 58862 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_15
timestamp 1607639953
transform 1 0 2466 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_3
timestamp 1607639953
transform 1 0 1362 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1607639953
transform 1 0 1086 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_39
timestamp 1607639953
transform 1 0 4674 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_27
timestamp 1607639953
transform 1 0 3570 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_62
timestamp 1607639953
transform 1 0 6790 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_59
timestamp 1607639953
transform 1 0 6514 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_89_51
timestamp 1607639953
transform 1 0 5778 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1104
timestamp 1607639953
transform 1 0 6698 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_86
timestamp 1607639953
transform 1 0 8998 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_74
timestamp 1607639953
transform 1 0 7894 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_110
timestamp 1607639953
transform 1 0 11206 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_98
timestamp 1607639953
transform 1 0 10102 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_123
timestamp 1607639953
transform 1 0 12402 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1105
timestamp 1607639953
transform 1 0 12310 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_147
timestamp 1607639953
transform 1 0 14610 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_135
timestamp 1607639953
transform 1 0 13506 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_171
timestamp 1607639953
transform 1 0 16818 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_159
timestamp 1607639953
transform 1 0 15714 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_187
timestamp 1607639953
transform 1 0 18290 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1106
timestamp 1607639953
transform 1 0 17922 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _106_
timestamp 1607639953
transform 1 0 18014 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_211
timestamp 1607639953
transform 1 0 20498 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_199
timestamp 1607639953
transform 1 0 19394 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_235
timestamp 1607639953
transform 1 0 22706 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_223
timestamp 1607639953
transform 1 0 21602 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_257
timestamp 1607639953
transform 1 0 24730 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_245
timestamp 1607639953
transform 1 0 23626 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_243
timestamp 1607639953
transform 1 0 23442 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1107
timestamp 1607639953
transform 1 0 23534 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_281
timestamp 1607639953
transform 1 0 26938 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_269
timestamp 1607639953
transform 1 0 25834 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_306
timestamp 1607639953
transform 1 0 29238 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_303
timestamp 1607639953
transform 1 0 28962 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_89_299
timestamp 1607639953
transform 1 0 28594 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_89_293
timestamp 1607639953
transform 1 0 28042 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1108
timestamp 1607639953
transform 1 0 29146 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _109_
timestamp 1607639953
transform 1 0 28686 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_330
timestamp 1607639953
transform 1 0 31446 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_318
timestamp 1607639953
transform 1 0 30342 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_342
timestamp 1607639953
transform 1 0 32550 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_367
timestamp 1607639953
transform 1 0 34850 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_354
timestamp 1607639953
transform 1 0 33654 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1109
timestamp 1607639953
transform 1 0 34758 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_391
timestamp 1607639953
transform 1 0 37058 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_379
timestamp 1607639953
transform 1 0 35954 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_415
timestamp 1607639953
transform 1 0 39266 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_403
timestamp 1607639953
transform 1 0 38162 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_440
timestamp 1607639953
transform 1 0 41566 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_428
timestamp 1607639953
transform 1 0 40462 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1110
timestamp 1607639953
transform 1 0 40370 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_452
timestamp 1607639953
transform 1 0 42670 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_476
timestamp 1607639953
transform 1 0 44878 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_464
timestamp 1607639953
transform 1 0 43774 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_501
timestamp 1607639953
transform 1 0 47178 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_489
timestamp 1607639953
transform 1 0 46074 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1111
timestamp 1607639953
transform 1 0 45982 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_525
timestamp 1607639953
transform 1 0 49386 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_513
timestamp 1607639953
transform 1 0 48282 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_550
timestamp 1607639953
transform 1 0 51686 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_537
timestamp 1607639953
transform 1 0 50490 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1112
timestamp 1607639953
transform 1 0 51594 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_562
timestamp 1607639953
transform 1 0 52790 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_586
timestamp 1607639953
transform 1 0 54998 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_574
timestamp 1607639953
transform 1 0 53894 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_611
timestamp 1607639953
transform 1 0 57298 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_598
timestamp 1607639953
transform 1 0 56102 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1113
timestamp 1607639953
transform 1 0 57206 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_623
timestamp 1607639953
transform 1 0 58402 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1607639953
transform -1 0 58862 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_15
timestamp 1607639953
transform 1 0 2466 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_3
timestamp 1607639953
transform 1 0 1362 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1607639953
transform 1 0 1086 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_44
timestamp 1607639953
transform 1 0 5134 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_32
timestamp 1607639953
transform 1 0 4030 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_27
timestamp 1607639953
transform 1 0 3570 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1114
timestamp 1607639953
transform 1 0 3938 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_56
timestamp 1607639953
transform 1 0 6238 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_80
timestamp 1607639953
transform 1 0 8446 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_68
timestamp 1607639953
transform 1 0 7342 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_107
timestamp 1607639953
transform 1 0 10930 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_90_101
timestamp 1607639953
transform 1 0 10378 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_90_93
timestamp 1607639953
transform 1 0 9642 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1115
timestamp 1607639953
transform 1 0 9550 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1607639953
transform 1 0 10654 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_131
timestamp 1607639953
transform 1 0 13138 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_119
timestamp 1607639953
transform 1 0 12034 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_154
timestamp 1607639953
transform 1 0 15254 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_151
timestamp 1607639953
transform 1 0 14978 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_90_143
timestamp 1607639953
transform 1 0 14242 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1116
timestamp 1607639953
transform 1 0 15162 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_166
timestamp 1607639953
transform 1 0 16358 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_190
timestamp 1607639953
transform 1 0 18566 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_178
timestamp 1607639953
transform 1 0 17462 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_215
timestamp 1607639953
transform 1 0 20866 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_202
timestamp 1607639953
transform 1 0 19670 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1117
timestamp 1607639953
transform 1 0 20774 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_239
timestamp 1607639953
transform 1 0 23074 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_227
timestamp 1607639953
transform 1 0 21970 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_263
timestamp 1607639953
transform 1 0 25282 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_251
timestamp 1607639953
transform 1 0 24178 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_276
timestamp 1607639953
transform 1 0 26478 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1118
timestamp 1607639953
transform 1 0 26386 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_300
timestamp 1607639953
transform 1 0 28686 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_288
timestamp 1607639953
transform 1 0 27582 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_324
timestamp 1607639953
transform 1 0 30894 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_312
timestamp 1607639953
transform 1 0 29790 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_349
timestamp 1607639953
transform 1 0 33194 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_337
timestamp 1607639953
transform 1 0 32090 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1119
timestamp 1607639953
transform 1 0 31998 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_373
timestamp 1607639953
transform 1 0 35402 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_361
timestamp 1607639953
transform 1 0 34298 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_385
timestamp 1607639953
transform 1 0 36506 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_410
timestamp 1607639953
transform 1 0 38806 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_398
timestamp 1607639953
transform 1 0 37702 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1120
timestamp 1607639953
transform 1 0 37610 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_434
timestamp 1607639953
transform 1 0 41014 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_422
timestamp 1607639953
transform 1 0 39910 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_459
timestamp 1607639953
transform 1 0 43314 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_446
timestamp 1607639953
transform 1 0 42118 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1121
timestamp 1607639953
transform 1 0 43222 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_483
timestamp 1607639953
transform 1 0 45522 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_471
timestamp 1607639953
transform 1 0 44418 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_495
timestamp 1607639953
transform 1 0 46626 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_520
timestamp 1607639953
transform 1 0 48926 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_507
timestamp 1607639953
transform 1 0 47730 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1122
timestamp 1607639953
transform 1 0 48834 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_544
timestamp 1607639953
transform 1 0 51134 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_532
timestamp 1607639953
transform 1 0 50030 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_568
timestamp 1607639953
transform 1 0 53342 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_556
timestamp 1607639953
transform 1 0 52238 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_593
timestamp 1607639953
transform 1 0 55642 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_581
timestamp 1607639953
transform 1 0 54538 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1123
timestamp 1607639953
transform 1 0 54446 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_605
timestamp 1607639953
transform 1 0 56746 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_617
timestamp 1607639953
transform 1 0 57850 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1607639953
transform -1 0 58862 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_15
timestamp 1607639953
transform 1 0 2466 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_3
timestamp 1607639953
transform 1 0 1362 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1607639953
transform 1 0 1086 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_39
timestamp 1607639953
transform 1 0 4674 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_27
timestamp 1607639953
transform 1 0 3570 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_62
timestamp 1607639953
transform 1 0 6790 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_59
timestamp 1607639953
transform 1 0 6514 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_91_51
timestamp 1607639953
transform 1 0 5778 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1124
timestamp 1607639953
transform 1 0 6698 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_86
timestamp 1607639953
transform 1 0 8998 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_74
timestamp 1607639953
transform 1 0 7894 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_110
timestamp 1607639953
transform 1 0 11206 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_98
timestamp 1607639953
transform 1 0 10102 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_123
timestamp 1607639953
transform 1 0 12402 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1125
timestamp 1607639953
transform 1 0 12310 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_147
timestamp 1607639953
transform 1 0 14610 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_135
timestamp 1607639953
transform 1 0 13506 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_171
timestamp 1607639953
transform 1 0 16818 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_159
timestamp 1607639953
transform 1 0 15714 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_196
timestamp 1607639953
transform 1 0 19118 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_184
timestamp 1607639953
transform 1 0 18014 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1126
timestamp 1607639953
transform 1 0 17922 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_220
timestamp 1607639953
transform 1 0 21326 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_208
timestamp 1607639953
transform 1 0 20222 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_232
timestamp 1607639953
transform 1 0 22430 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_257
timestamp 1607639953
transform 1 0 24730 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_245
timestamp 1607639953
transform 1 0 23626 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1127
timestamp 1607639953
transform 1 0 23534 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_281
timestamp 1607639953
transform 1 0 26938 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_269
timestamp 1607639953
transform 1 0 25834 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_306
timestamp 1607639953
transform 1 0 29238 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_293
timestamp 1607639953
transform 1 0 28042 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1128
timestamp 1607639953
transform 1 0 29146 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_330
timestamp 1607639953
transform 1 0 31446 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_318
timestamp 1607639953
transform 1 0 30342 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_342
timestamp 1607639953
transform 1 0 32550 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_367
timestamp 1607639953
transform 1 0 34850 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_354
timestamp 1607639953
transform 1 0 33654 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1129
timestamp 1607639953
transform 1 0 34758 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_391
timestamp 1607639953
transform 1 0 37058 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_379
timestamp 1607639953
transform 1 0 35954 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_415
timestamp 1607639953
transform 1 0 39266 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_403
timestamp 1607639953
transform 1 0 38162 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_440
timestamp 1607639953
transform 1 0 41566 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_428
timestamp 1607639953
transform 1 0 40462 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1130
timestamp 1607639953
transform 1 0 40370 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_452
timestamp 1607639953
transform 1 0 42670 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_476
timestamp 1607639953
transform 1 0 44878 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_464
timestamp 1607639953
transform 1 0 43774 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_501
timestamp 1607639953
transform 1 0 47178 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_489
timestamp 1607639953
transform 1 0 46074 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1131
timestamp 1607639953
transform 1 0 45982 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_525
timestamp 1607639953
transform 1 0 49386 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_513
timestamp 1607639953
transform 1 0 48282 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_550
timestamp 1607639953
transform 1 0 51686 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_537
timestamp 1607639953
transform 1 0 50490 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1132
timestamp 1607639953
transform 1 0 51594 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_562
timestamp 1607639953
transform 1 0 52790 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_586
timestamp 1607639953
transform 1 0 54998 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_574
timestamp 1607639953
transform 1 0 53894 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_611
timestamp 1607639953
transform 1 0 57298 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_598
timestamp 1607639953
transform 1 0 56102 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1133
timestamp 1607639953
transform 1 0 57206 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_623
timestamp 1607639953
transform 1 0 58402 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1607639953
transform -1 0 58862 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_15
timestamp 1607639953
transform 1 0 2466 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_3
timestamp 1607639953
transform 1 0 1362 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_15
timestamp 1607639953
transform 1 0 2466 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_3
timestamp 1607639953
transform 1 0 1362 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1607639953
transform 1 0 1086 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1607639953
transform 1 0 1086 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_39
timestamp 1607639953
transform 1 0 4674 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_27
timestamp 1607639953
transform 1 0 3570 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_44
timestamp 1607639953
transform 1 0 5134 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_32
timestamp 1607639953
transform 1 0 4030 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_27
timestamp 1607639953
transform 1 0 3570 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1134
timestamp 1607639953
transform 1 0 3938 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_62
timestamp 1607639953
transform 1 0 6790 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_59
timestamp 1607639953
transform 1 0 6514 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_51
timestamp 1607639953
transform 1 0 5778 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_56
timestamp 1607639953
transform 1 0 6238 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1144
timestamp 1607639953
transform 1 0 6698 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_86
timestamp 1607639953
transform 1 0 8998 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_74
timestamp 1607639953
transform 1 0 7894 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_84
timestamp 1607639953
transform 1 0 8814 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_72
timestamp 1607639953
transform 1 0 7710 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_68
timestamp 1607639953
transform 1 0 7342 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _128_
timestamp 1607639953
transform 1 0 7434 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_110
timestamp 1607639953
transform 1 0 11206 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_98
timestamp 1607639953
transform 1 0 10102 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_105
timestamp 1607639953
transform 1 0 10746 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_93
timestamp 1607639953
transform 1 0 9642 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1135
timestamp 1607639953
transform 1 0 9550 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_123
timestamp 1607639953
transform 1 0 12402 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_131
timestamp 1607639953
transform 1 0 13138 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_119
timestamp 1607639953
transform 1 0 12034 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_92_113
timestamp 1607639953
transform 1 0 11482 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1145
timestamp 1607639953
transform 1 0 12310 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _185_
timestamp 1607639953
transform 1 0 11758 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_153
timestamp 1607639953
transform 1 0 15162 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_141
timestamp 1607639953
transform 1 0 14058 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_135
timestamp 1607639953
transform 1 0 13506 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_154
timestamp 1607639953
transform 1 0 15254 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_151
timestamp 1607639953
transform 1 0 14978 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_92_143
timestamp 1607639953
transform 1 0 14242 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1136
timestamp 1607639953
transform 1 0 15162 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _202_
timestamp 1607639953
transform 1 0 13782 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_165
timestamp 1607639953
transform 1 0 16266 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_166
timestamp 1607639953
transform 1 0 16358 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_190
timestamp 1607639953
transform 1 0 18566 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_184
timestamp 1607639953
transform 1 0 18014 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_93_177
timestamp 1607639953
transform 1 0 17370 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_92_190
timestamp 1607639953
transform 1 0 18566 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_178
timestamp 1607639953
transform 1 0 17462 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1146
timestamp 1607639953
transform 1 0 17922 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _027_
timestamp 1607639953
transform 1 0 18290 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_214
timestamp 1607639953
transform 1 0 20774 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_202
timestamp 1607639953
transform 1 0 19670 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_215
timestamp 1607639953
transform 1 0 20866 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_202
timestamp 1607639953
transform 1 0 19670 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1137
timestamp 1607639953
transform 1 0 20774 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_93_238
timestamp 1607639953
transform 1 0 22982 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_93_226
timestamp 1607639953
transform 1 0 21878 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_239
timestamp 1607639953
transform 1 0 23074 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_227
timestamp 1607639953
transform 1 0 21970 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_257
timestamp 1607639953
transform 1 0 24730 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_245
timestamp 1607639953
transform 1 0 23626 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_263
timestamp 1607639953
transform 1 0 25282 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_251
timestamp 1607639953
transform 1 0 24178 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1147
timestamp 1607639953
transform 1 0 23534 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_281
timestamp 1607639953
transform 1 0 26938 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_269
timestamp 1607639953
transform 1 0 25834 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_276
timestamp 1607639953
transform 1 0 26478 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1138
timestamp 1607639953
transform 1 0 26386 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_306
timestamp 1607639953
transform 1 0 29238 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_293
timestamp 1607639953
transform 1 0 28042 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_300
timestamp 1607639953
transform 1 0 28686 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_288
timestamp 1607639953
transform 1 0 27582 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1148
timestamp 1607639953
transform 1 0 29146 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_330
timestamp 1607639953
transform 1 0 31446 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_318
timestamp 1607639953
transform 1 0 30342 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_324
timestamp 1607639953
transform 1 0 30894 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_312
timestamp 1607639953
transform 1 0 29790 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_342
timestamp 1607639953
transform 1 0 32550 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_349
timestamp 1607639953
transform 1 0 33194 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_345
timestamp 1607639953
transform 1 0 32826 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_337
timestamp 1607639953
transform 1 0 32090 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1139
timestamp 1607639953
transform 1 0 31998 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1607639953
transform 1 0 32918 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_367
timestamp 1607639953
transform 1 0 34850 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_354
timestamp 1607639953
transform 1 0 33654 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_373
timestamp 1607639953
transform 1 0 35402 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_361
timestamp 1607639953
transform 1 0 34298 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1149
timestamp 1607639953
transform 1 0 34758 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_391
timestamp 1607639953
transform 1 0 37058 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_379
timestamp 1607639953
transform 1 0 35954 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_385
timestamp 1607639953
transform 1 0 36506 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_415
timestamp 1607639953
transform 1 0 39266 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_403
timestamp 1607639953
transform 1 0 38162 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_416
timestamp 1607639953
transform 1 0 39358 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_410
timestamp 1607639953
transform 1 0 38806 0 -1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_92_398
timestamp 1607639953
transform 1 0 37702 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1140
timestamp 1607639953
transform 1 0 37610 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _155_
timestamp 1607639953
transform 1 0 39450 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_440
timestamp 1607639953
transform 1 0 41566 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_428
timestamp 1607639953
transform 1 0 40462 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_432
timestamp 1607639953
transform 1 0 40830 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_420
timestamp 1607639953
transform 1 0 39726 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1150
timestamp 1607639953
transform 1 0 40370 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_452
timestamp 1607639953
transform 1 0 42670 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_459
timestamp 1607639953
transform 1 0 43314 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_456
timestamp 1607639953
transform 1 0 43038 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_92_444
timestamp 1607639953
transform 1 0 41934 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1141
timestamp 1607639953
transform 1 0 43222 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_476
timestamp 1607639953
transform 1 0 44878 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_464
timestamp 1607639953
transform 1 0 43774 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_483
timestamp 1607639953
transform 1 0 45522 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_471
timestamp 1607639953
transform 1 0 44418 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_501
timestamp 1607639953
transform 1 0 47178 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_489
timestamp 1607639953
transform 1 0 46074 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_495
timestamp 1607639953
transform 1 0 46626 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1151
timestamp 1607639953
transform 1 0 45982 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_525
timestamp 1607639953
transform 1 0 49386 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_513
timestamp 1607639953
transform 1 0 48282 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_520
timestamp 1607639953
transform 1 0 48926 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_507
timestamp 1607639953
transform 1 0 47730 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1142
timestamp 1607639953
transform 1 0 48834 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_550
timestamp 1607639953
transform 1 0 51686 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_537
timestamp 1607639953
transform 1 0 50490 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_544
timestamp 1607639953
transform 1 0 51134 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_532
timestamp 1607639953
transform 1 0 50030 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1152
timestamp 1607639953
transform 1 0 51594 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_562
timestamp 1607639953
transform 1 0 52790 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_568
timestamp 1607639953
transform 1 0 53342 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_556
timestamp 1607639953
transform 1 0 52238 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_586
timestamp 1607639953
transform 1 0 54998 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_574
timestamp 1607639953
transform 1 0 53894 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_593
timestamp 1607639953
transform 1 0 55642 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_581
timestamp 1607639953
transform 1 0 54538 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1143
timestamp 1607639953
transform 1 0 54446 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_611
timestamp 1607639953
transform 1 0 57298 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_598
timestamp 1607639953
transform 1 0 56102 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_605
timestamp 1607639953
transform 1 0 56746 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1153
timestamp 1607639953
transform 1 0 57206 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_623
timestamp 1607639953
transform 1 0 58402 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_92_617
timestamp 1607639953
transform 1 0 57850 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1607639953
transform -1 0 58862 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1607639953
transform -1 0 58862 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_15
timestamp 1607639953
transform 1 0 2466 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_3
timestamp 1607639953
transform 1 0 1362 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1607639953
transform 1 0 1086 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_44
timestamp 1607639953
transform 1 0 5134 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_32
timestamp 1607639953
transform 1 0 4030 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_27
timestamp 1607639953
transform 1 0 3570 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1154
timestamp 1607639953
transform 1 0 3938 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_56
timestamp 1607639953
transform 1 0 6238 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_80
timestamp 1607639953
transform 1 0 8446 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_68
timestamp 1607639953
transform 1 0 7342 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_105
timestamp 1607639953
transform 1 0 10746 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_93
timestamp 1607639953
transform 1 0 9642 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1155
timestamp 1607639953
transform 1 0 9550 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_129
timestamp 1607639953
transform 1 0 12954 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_117
timestamp 1607639953
transform 1 0 11850 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_154
timestamp 1607639953
transform 1 0 15254 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_141
timestamp 1607639953
transform 1 0 14058 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1156
timestamp 1607639953
transform 1 0 15162 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_166
timestamp 1607639953
transform 1 0 16358 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_190
timestamp 1607639953
transform 1 0 18566 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_178
timestamp 1607639953
transform 1 0 17462 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_215
timestamp 1607639953
transform 1 0 20866 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_202
timestamp 1607639953
transform 1 0 19670 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1157
timestamp 1607639953
transform 1 0 20774 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_94_239
timestamp 1607639953
transform 1 0 23074 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_94_227
timestamp 1607639953
transform 1 0 21970 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_260
timestamp 1607639953
transform 1 0 25006 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_248
timestamp 1607639953
transform 1 0 23902 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _004_
timestamp 1607639953
transform 1 0 23626 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_276
timestamp 1607639953
transform 1 0 26478 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_94_272
timestamp 1607639953
transform 1 0 26110 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1158
timestamp 1607639953
transform 1 0 26386 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_300
timestamp 1607639953
transform 1 0 28686 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_288
timestamp 1607639953
transform 1 0 27582 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_324
timestamp 1607639953
transform 1 0 30894 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_312
timestamp 1607639953
transform 1 0 29790 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_349
timestamp 1607639953
transform 1 0 33194 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_337
timestamp 1607639953
transform 1 0 32090 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1159
timestamp 1607639953
transform 1 0 31998 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_373
timestamp 1607639953
transform 1 0 35402 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_361
timestamp 1607639953
transform 1 0 34298 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_385
timestamp 1607639953
transform 1 0 36506 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_410
timestamp 1607639953
transform 1 0 38806 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_398
timestamp 1607639953
transform 1 0 37702 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1160
timestamp 1607639953
transform 1 0 37610 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_434
timestamp 1607639953
transform 1 0 41014 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_422
timestamp 1607639953
transform 1 0 39910 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_459
timestamp 1607639953
transform 1 0 43314 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_446
timestamp 1607639953
transform 1 0 42118 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1161
timestamp 1607639953
transform 1 0 43222 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_483
timestamp 1607639953
transform 1 0 45522 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_471
timestamp 1607639953
transform 1 0 44418 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_495
timestamp 1607639953
transform 1 0 46626 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_520
timestamp 1607639953
transform 1 0 48926 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_507
timestamp 1607639953
transform 1 0 47730 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1162
timestamp 1607639953
transform 1 0 48834 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_544
timestamp 1607639953
transform 1 0 51134 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_532
timestamp 1607639953
transform 1 0 50030 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_568
timestamp 1607639953
transform 1 0 53342 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_556
timestamp 1607639953
transform 1 0 52238 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_593
timestamp 1607639953
transform 1 0 55642 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_581
timestamp 1607639953
transform 1 0 54538 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1163
timestamp 1607639953
transform 1 0 54446 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_605
timestamp 1607639953
transform 1 0 56746 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_617
timestamp 1607639953
transform 1 0 57850 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1607639953
transform -1 0 58862 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_18
timestamp 1607639953
transform 1 0 2742 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_6
timestamp 1607639953
transform 1 0 1638 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1607639953
transform 1 0 1086 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _085_
timestamp 1607639953
transform 1 0 1362 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_42
timestamp 1607639953
transform 1 0 4950 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_30
timestamp 1607639953
transform 1 0 3846 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_62
timestamp 1607639953
transform 1 0 6790 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_95_60
timestamp 1607639953
transform 1 0 6606 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_95_54
timestamp 1607639953
transform 1 0 6054 0 1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1164
timestamp 1607639953
transform 1 0 6698 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_86
timestamp 1607639953
transform 1 0 8998 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_74
timestamp 1607639953
transform 1 0 7894 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_110
timestamp 1607639953
transform 1 0 11206 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_98
timestamp 1607639953
transform 1 0 10102 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_123
timestamp 1607639953
transform 1 0 12402 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1165
timestamp 1607639953
transform 1 0 12310 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_147
timestamp 1607639953
transform 1 0 14610 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_135
timestamp 1607639953
transform 1 0 13506 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_171
timestamp 1607639953
transform 1 0 16818 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_159
timestamp 1607639953
transform 1 0 15714 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_196
timestamp 1607639953
transform 1 0 19118 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_184
timestamp 1607639953
transform 1 0 18014 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1166
timestamp 1607639953
transform 1 0 17922 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_220
timestamp 1607639953
transform 1 0 21326 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_208
timestamp 1607639953
transform 1 0 20222 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_232
timestamp 1607639953
transform 1 0 22430 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_257
timestamp 1607639953
transform 1 0 24730 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_245
timestamp 1607639953
transform 1 0 23626 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1167
timestamp 1607639953
transform 1 0 23534 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_281
timestamp 1607639953
transform 1 0 26938 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_269
timestamp 1607639953
transform 1 0 25834 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_306
timestamp 1607639953
transform 1 0 29238 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_293
timestamp 1607639953
transform 1 0 28042 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1168
timestamp 1607639953
transform 1 0 29146 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_330
timestamp 1607639953
transform 1 0 31446 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_318
timestamp 1607639953
transform 1 0 30342 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_342
timestamp 1607639953
transform 1 0 32550 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_367
timestamp 1607639953
transform 1 0 34850 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_354
timestamp 1607639953
transform 1 0 33654 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1169
timestamp 1607639953
transform 1 0 34758 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_391
timestamp 1607639953
transform 1 0 37058 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_379
timestamp 1607639953
transform 1 0 35954 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_415
timestamp 1607639953
transform 1 0 39266 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_403
timestamp 1607639953
transform 1 0 38162 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_440
timestamp 1607639953
transform 1 0 41566 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_428
timestamp 1607639953
transform 1 0 40462 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1170
timestamp 1607639953
transform 1 0 40370 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_452
timestamp 1607639953
transform 1 0 42670 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_476
timestamp 1607639953
transform 1 0 44878 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_464
timestamp 1607639953
transform 1 0 43774 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_501
timestamp 1607639953
transform 1 0 47178 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_489
timestamp 1607639953
transform 1 0 46074 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1171
timestamp 1607639953
transform 1 0 45982 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_525
timestamp 1607639953
transform 1 0 49386 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_513
timestamp 1607639953
transform 1 0 48282 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_550
timestamp 1607639953
transform 1 0 51686 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_537
timestamp 1607639953
transform 1 0 50490 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1172
timestamp 1607639953
transform 1 0 51594 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_562
timestamp 1607639953
transform 1 0 52790 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_586
timestamp 1607639953
transform 1 0 54998 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_574
timestamp 1607639953
transform 1 0 53894 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_611
timestamp 1607639953
transform 1 0 57298 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_598
timestamp 1607639953
transform 1 0 56102 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1173
timestamp 1607639953
transform 1 0 57206 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_623
timestamp 1607639953
transform 1 0 58402 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1607639953
transform -1 0 58862 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_15
timestamp 1607639953
transform 1 0 2466 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_3
timestamp 1607639953
transform 1 0 1362 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1607639953
transform 1 0 1086 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_44
timestamp 1607639953
transform 1 0 5134 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_32
timestamp 1607639953
transform 1 0 4030 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_27
timestamp 1607639953
transform 1 0 3570 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1174
timestamp 1607639953
transform 1 0 3938 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_56
timestamp 1607639953
transform 1 0 6238 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_80
timestamp 1607639953
transform 1 0 8446 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_68
timestamp 1607639953
transform 1 0 7342 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_105
timestamp 1607639953
transform 1 0 10746 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_93
timestamp 1607639953
transform 1 0 9642 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1175
timestamp 1607639953
transform 1 0 9550 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_129
timestamp 1607639953
transform 1 0 12954 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_117
timestamp 1607639953
transform 1 0 11850 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_154
timestamp 1607639953
transform 1 0 15254 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_141
timestamp 1607639953
transform 1 0 14058 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1176
timestamp 1607639953
transform 1 0 15162 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_166
timestamp 1607639953
transform 1 0 16358 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_198
timestamp 1607639953
transform 1 0 19302 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_186
timestamp 1607639953
transform 1 0 18198 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_182
timestamp 1607639953
transform 1 0 17830 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_178
timestamp 1607639953
transform 1 0 17462 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _112_
timestamp 1607639953
transform 1 0 17922 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_218
timestamp 1607639953
transform 1 0 21142 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_210
timestamp 1607639953
transform 1 0 20406 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1177
timestamp 1607639953
transform 1 0 20774 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _164_
timestamp 1607639953
transform 1 0 20866 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_242
timestamp 1607639953
transform 1 0 23350 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_230
timestamp 1607639953
transform 1 0 22246 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_254
timestamp 1607639953
transform 1 0 24454 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_276
timestamp 1607639953
transform 1 0 26478 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_274
timestamp 1607639953
transform 1 0 26294 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_266
timestamp 1607639953
transform 1 0 25558 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1178
timestamp 1607639953
transform 1 0 26386 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_300
timestamp 1607639953
transform 1 0 28686 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_288
timestamp 1607639953
transform 1 0 27582 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_324
timestamp 1607639953
transform 1 0 30894 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_312
timestamp 1607639953
transform 1 0 29790 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_349
timestamp 1607639953
transform 1 0 33194 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_337
timestamp 1607639953
transform 1 0 32090 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1179
timestamp 1607639953
transform 1 0 31998 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_373
timestamp 1607639953
transform 1 0 35402 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_361
timestamp 1607639953
transform 1 0 34298 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_385
timestamp 1607639953
transform 1 0 36506 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_410
timestamp 1607639953
transform 1 0 38806 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_398
timestamp 1607639953
transform 1 0 37702 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1180
timestamp 1607639953
transform 1 0 37610 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_434
timestamp 1607639953
transform 1 0 41014 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_422
timestamp 1607639953
transform 1 0 39910 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_96_459
timestamp 1607639953
transform 1 0 43314 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_446
timestamp 1607639953
transform 1 0 42118 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1181
timestamp 1607639953
transform 1 0 43222 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _179_
timestamp 1607639953
transform 1 0 43590 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_477
timestamp 1607639953
transform 1 0 44970 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_465
timestamp 1607639953
transform 1 0 43866 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_501
timestamp 1607639953
transform 1 0 47178 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_489
timestamp 1607639953
transform 1 0 46074 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_520
timestamp 1607639953
transform 1 0 48926 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_513
timestamp 1607639953
transform 1 0 48282 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1182
timestamp 1607639953
transform 1 0 48834 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_544
timestamp 1607639953
transform 1 0 51134 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_532
timestamp 1607639953
transform 1 0 50030 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_568
timestamp 1607639953
transform 1 0 53342 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_556
timestamp 1607639953
transform 1 0 52238 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_593
timestamp 1607639953
transform 1 0 55642 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_581
timestamp 1607639953
transform 1 0 54538 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1183
timestamp 1607639953
transform 1 0 54446 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_605
timestamp 1607639953
transform 1 0 56746 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_617
timestamp 1607639953
transform 1 0 57850 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1607639953
transform -1 0 58862 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_15
timestamp 1607639953
transform 1 0 2466 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_3
timestamp 1607639953
transform 1 0 1362 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1607639953
transform 1 0 1086 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_39
timestamp 1607639953
transform 1 0 4674 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_27
timestamp 1607639953
transform 1 0 3570 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_62
timestamp 1607639953
transform 1 0 6790 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_59
timestamp 1607639953
transform 1 0 6514 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_97_51
timestamp 1607639953
transform 1 0 5778 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1184
timestamp 1607639953
transform 1 0 6698 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_86
timestamp 1607639953
transform 1 0 8998 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_74
timestamp 1607639953
transform 1 0 7894 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_110
timestamp 1607639953
transform 1 0 11206 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_98
timestamp 1607639953
transform 1 0 10102 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_123
timestamp 1607639953
transform 1 0 12402 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1185
timestamp 1607639953
transform 1 0 12310 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_147
timestamp 1607639953
transform 1 0 14610 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_135
timestamp 1607639953
transform 1 0 13506 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_171
timestamp 1607639953
transform 1 0 16818 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_159
timestamp 1607639953
transform 1 0 15714 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_196
timestamp 1607639953
transform 1 0 19118 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_184
timestamp 1607639953
transform 1 0 18014 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1186
timestamp 1607639953
transform 1 0 17922 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_220
timestamp 1607639953
transform 1 0 21326 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_208
timestamp 1607639953
transform 1 0 20222 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_232
timestamp 1607639953
transform 1 0 22430 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_257
timestamp 1607639953
transform 1 0 24730 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_245
timestamp 1607639953
transform 1 0 23626 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1187
timestamp 1607639953
transform 1 0 23534 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_281
timestamp 1607639953
transform 1 0 26938 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_269
timestamp 1607639953
transform 1 0 25834 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_306
timestamp 1607639953
transform 1 0 29238 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_293
timestamp 1607639953
transform 1 0 28042 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1188
timestamp 1607639953
transform 1 0 29146 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_330
timestamp 1607639953
transform 1 0 31446 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_318
timestamp 1607639953
transform 1 0 30342 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_342
timestamp 1607639953
transform 1 0 32550 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_367
timestamp 1607639953
transform 1 0 34850 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_354
timestamp 1607639953
transform 1 0 33654 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1189
timestamp 1607639953
transform 1 0 34758 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_391
timestamp 1607639953
transform 1 0 37058 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_379
timestamp 1607639953
transform 1 0 35954 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_415
timestamp 1607639953
transform 1 0 39266 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_403
timestamp 1607639953
transform 1 0 38162 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_440
timestamp 1607639953
transform 1 0 41566 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_428
timestamp 1607639953
transform 1 0 40462 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1190
timestamp 1607639953
transform 1 0 40370 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_452
timestamp 1607639953
transform 1 0 42670 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_476
timestamp 1607639953
transform 1 0 44878 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_464
timestamp 1607639953
transform 1 0 43774 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_501
timestamp 1607639953
transform 1 0 47178 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_489
timestamp 1607639953
transform 1 0 46074 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1191
timestamp 1607639953
transform 1 0 45982 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_525
timestamp 1607639953
transform 1 0 49386 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_513
timestamp 1607639953
transform 1 0 48282 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_550
timestamp 1607639953
transform 1 0 51686 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_537
timestamp 1607639953
transform 1 0 50490 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1192
timestamp 1607639953
transform 1 0 51594 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_562
timestamp 1607639953
transform 1 0 52790 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_586
timestamp 1607639953
transform 1 0 54998 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_574
timestamp 1607639953
transform 1 0 53894 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_611
timestamp 1607639953
transform 1 0 57298 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_598
timestamp 1607639953
transform 1 0 56102 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1193
timestamp 1607639953
transform 1 0 57206 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_623
timestamp 1607639953
transform 1 0 58402 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1607639953
transform -1 0 58862 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_15
timestamp 1607639953
transform 1 0 2466 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_3
timestamp 1607639953
transform 1 0 1362 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1607639953
transform 1 0 1086 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_44
timestamp 1607639953
transform 1 0 5134 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_32
timestamp 1607639953
transform 1 0 4030 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_27
timestamp 1607639953
transform 1 0 3570 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1194
timestamp 1607639953
transform 1 0 3938 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_56
timestamp 1607639953
transform 1 0 6238 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_80
timestamp 1607639953
transform 1 0 8446 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_68
timestamp 1607639953
transform 1 0 7342 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_105
timestamp 1607639953
transform 1 0 10746 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_93
timestamp 1607639953
transform 1 0 9642 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1195
timestamp 1607639953
transform 1 0 9550 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_129
timestamp 1607639953
transform 1 0 12954 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_117
timestamp 1607639953
transform 1 0 11850 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_154
timestamp 1607639953
transform 1 0 15254 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_141
timestamp 1607639953
transform 1 0 14058 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1196
timestamp 1607639953
transform 1 0 15162 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_166
timestamp 1607639953
transform 1 0 16358 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_190
timestamp 1607639953
transform 1 0 18566 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_178
timestamp 1607639953
transform 1 0 17462 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_215
timestamp 1607639953
transform 1 0 20866 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_202
timestamp 1607639953
transform 1 0 19670 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1197
timestamp 1607639953
transform 1 0 20774 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_239
timestamp 1607639953
transform 1 0 23074 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_227
timestamp 1607639953
transform 1 0 21970 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_263
timestamp 1607639953
transform 1 0 25282 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_251
timestamp 1607639953
transform 1 0 24178 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_276
timestamp 1607639953
transform 1 0 26478 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1198
timestamp 1607639953
transform 1 0 26386 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_305
timestamp 1607639953
transform 1 0 29146 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_293
timestamp 1607639953
transform 1 0 28042 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_98_288
timestamp 1607639953
transform 1 0 27582 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1607639953
transform 1 0 27766 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_98_329
timestamp 1607639953
transform 1 0 31354 0 -1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_98_317
timestamp 1607639953
transform 1 0 30250 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_349
timestamp 1607639953
transform 1 0 33194 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_337
timestamp 1607639953
transform 1 0 32090 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_335
timestamp 1607639953
transform 1 0 31906 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1199
timestamp 1607639953
transform 1 0 31998 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_373
timestamp 1607639953
transform 1 0 35402 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_361
timestamp 1607639953
transform 1 0 34298 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_385
timestamp 1607639953
transform 1 0 36506 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_413
timestamp 1607639953
transform 1 0 39082 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_401
timestamp 1607639953
transform 1 0 37978 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1200
timestamp 1607639953
transform 1 0 37610 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _024_
timestamp 1607639953
transform 1 0 37702 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_437
timestamp 1607639953
transform 1 0 41290 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_425
timestamp 1607639953
transform 1 0 40186 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_459
timestamp 1607639953
transform 1 0 43314 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_457
timestamp 1607639953
transform 1 0 43130 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_449
timestamp 1607639953
transform 1 0 42394 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1201
timestamp 1607639953
transform 1 0 43222 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_483
timestamp 1607639953
transform 1 0 45522 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_471
timestamp 1607639953
transform 1 0 44418 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_495
timestamp 1607639953
transform 1 0 46626 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_520
timestamp 1607639953
transform 1 0 48926 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_507
timestamp 1607639953
transform 1 0 47730 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1202
timestamp 1607639953
transform 1 0 48834 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_544
timestamp 1607639953
transform 1 0 51134 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_532
timestamp 1607639953
transform 1 0 50030 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_571
timestamp 1607639953
transform 1 0 53618 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_559
timestamp 1607639953
transform 1 0 52514 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _153_
timestamp 1607639953
transform 1 0 52238 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_593
timestamp 1607639953
transform 1 0 55642 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_581
timestamp 1607639953
transform 1 0 54538 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_579
timestamp 1607639953
transform 1 0 54354 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1203
timestamp 1607639953
transform 1 0 54446 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_605
timestamp 1607639953
transform 1 0 56746 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_617
timestamp 1607639953
transform 1 0 57850 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1607639953
transform -1 0 58862 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_18
timestamp 1607639953
transform 1 0 2742 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_3
timestamp 1607639953
transform 1 0 1362 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_15
timestamp 1607639953
transform 1 0 2466 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_3
timestamp 1607639953
transform 1 0 1362 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1607639953
transform 1 0 1086 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1607639953
transform 1 0 1086 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1607639953
transform 1 0 2466 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_44
timestamp 1607639953
transform 1 0 5134 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_32
timestamp 1607639953
transform 1 0 4030 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_30
timestamp 1607639953
transform 1 0 3846 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_39
timestamp 1607639953
transform 1 0 4674 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_27
timestamp 1607639953
transform 1 0 3570 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1214
timestamp 1607639953
transform 1 0 3938 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_56
timestamp 1607639953
transform 1 0 6238 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_62
timestamp 1607639953
transform 1 0 6790 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_58
timestamp 1607639953
transform 1 0 6422 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1607639953
transform 1 0 5778 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1204
timestamp 1607639953
transform 1 0 6698 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _008_
timestamp 1607639953
transform 1 0 6146 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_80
timestamp 1607639953
transform 1 0 8446 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_68
timestamp 1607639953
transform 1 0 7342 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_86
timestamp 1607639953
transform 1 0 8998 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_74
timestamp 1607639953
transform 1 0 7894 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_108
timestamp 1607639953
transform 1 0 11022 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_96
timestamp 1607639953
transform 1 0 9918 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_110
timestamp 1607639953
transform 1 0 11206 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_98
timestamp 1607639953
transform 1 0 10102 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1215
timestamp 1607639953
transform 1 0 9550 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _007_
timestamp 1607639953
transform 1 0 9642 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_132
timestamp 1607639953
transform 1 0 13230 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_120
timestamp 1607639953
transform 1 0 12126 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_123
timestamp 1607639953
transform 1 0 12402 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1205
timestamp 1607639953
transform 1 0 12310 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_154
timestamp 1607639953
transform 1 0 15254 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_152
timestamp 1607639953
transform 1 0 15070 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_144
timestamp 1607639953
transform 1 0 14334 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_147
timestamp 1607639953
transform 1 0 14610 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_135
timestamp 1607639953
transform 1 0 13506 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1216
timestamp 1607639953
transform 1 0 15162 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_166
timestamp 1607639953
transform 1 0 16358 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_169
timestamp 1607639953
transform 1 0 16634 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_165
timestamp 1607639953
transform 1 0 16266 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_99_159
timestamp 1607639953
transform 1 0 15714 0 1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _073_
timestamp 1607639953
transform 1 0 16358 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_190
timestamp 1607639953
transform 1 0 18566 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_178
timestamp 1607639953
transform 1 0 17462 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_196
timestamp 1607639953
transform 1 0 19118 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_184
timestamp 1607639953
transform 1 0 18014 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_181
timestamp 1607639953
transform 1 0 17738 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1206
timestamp 1607639953
transform 1 0 17922 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_215
timestamp 1607639953
transform 1 0 20866 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_202
timestamp 1607639953
transform 1 0 19670 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_220
timestamp 1607639953
transform 1 0 21326 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_208
timestamp 1607639953
transform 1 0 20222 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1217
timestamp 1607639953
transform 1 0 20774 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_239
timestamp 1607639953
transform 1 0 23074 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_227
timestamp 1607639953
transform 1 0 21970 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_232
timestamp 1607639953
transform 1 0 22430 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_263
timestamp 1607639953
transform 1 0 25282 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_251
timestamp 1607639953
transform 1 0 24178 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_257
timestamp 1607639953
transform 1 0 24730 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_245
timestamp 1607639953
transform 1 0 23626 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1207
timestamp 1607639953
transform 1 0 23534 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_276
timestamp 1607639953
transform 1 0 26478 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_281
timestamp 1607639953
transform 1 0 26938 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_269
timestamp 1607639953
transform 1 0 25834 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1218
timestamp 1607639953
transform 1 0 26386 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_300
timestamp 1607639953
transform 1 0 28686 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_288
timestamp 1607639953
transform 1 0 27582 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_306
timestamp 1607639953
transform 1 0 29238 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_293
timestamp 1607639953
transform 1 0 28042 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1208
timestamp 1607639953
transform 1 0 29146 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _020_
timestamp 1607639953
transform 1 0 29422 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_323
timestamp 1607639953
transform 1 0 30802 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_311
timestamp 1607639953
transform 1 0 29698 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_330
timestamp 1607639953
transform 1 0 31446 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_318
timestamp 1607639953
transform 1 0 30342 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_349
timestamp 1607639953
transform 1 0 33194 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_337
timestamp 1607639953
transform 1 0 32090 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_335
timestamp 1607639953
transform 1 0 31906 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_342
timestamp 1607639953
transform 1 0 32550 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1219
timestamp 1607639953
transform 1 0 31998 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_373
timestamp 1607639953
transform 1 0 35402 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_361
timestamp 1607639953
transform 1 0 34298 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_367
timestamp 1607639953
transform 1 0 34850 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_354
timestamp 1607639953
transform 1 0 33654 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1209
timestamp 1607639953
transform 1 0 34758 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_385
timestamp 1607639953
transform 1 0 36506 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_391
timestamp 1607639953
transform 1 0 37058 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_379
timestamp 1607639953
transform 1 0 35954 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_410
timestamp 1607639953
transform 1 0 38806 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_398
timestamp 1607639953
transform 1 0 37702 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_415
timestamp 1607639953
transform 1 0 39266 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_403
timestamp 1607639953
transform 1 0 38162 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1220
timestamp 1607639953
transform 1 0 37610 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_434
timestamp 1607639953
transform 1 0 41014 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_422
timestamp 1607639953
transform 1 0 39910 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_440
timestamp 1607639953
transform 1 0 41566 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_428
timestamp 1607639953
transform 1 0 40462 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1210
timestamp 1607639953
transform 1 0 40370 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_459
timestamp 1607639953
transform 1 0 43314 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_446
timestamp 1607639953
transform 1 0 42118 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_452
timestamp 1607639953
transform 1 0 42670 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1221
timestamp 1607639953
transform 1 0 43222 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_483
timestamp 1607639953
transform 1 0 45522 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_471
timestamp 1607639953
transform 1 0 44418 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_476
timestamp 1607639953
transform 1 0 44878 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_464
timestamp 1607639953
transform 1 0 43774 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_495
timestamp 1607639953
transform 1 0 46626 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_501
timestamp 1607639953
transform 1 0 47178 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_489
timestamp 1607639953
transform 1 0 46074 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1211
timestamp 1607639953
transform 1 0 45982 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_520
timestamp 1607639953
transform 1 0 48926 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_507
timestamp 1607639953
transform 1 0 47730 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_525
timestamp 1607639953
transform 1 0 49386 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_513
timestamp 1607639953
transform 1 0 48282 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1222
timestamp 1607639953
transform 1 0 48834 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_544
timestamp 1607639953
transform 1 0 51134 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_532
timestamp 1607639953
transform 1 0 50030 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_550
timestamp 1607639953
transform 1 0 51686 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_537
timestamp 1607639953
transform 1 0 50490 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1212
timestamp 1607639953
transform 1 0 51594 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_568
timestamp 1607639953
transform 1 0 53342 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_556
timestamp 1607639953
transform 1 0 52238 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_562
timestamp 1607639953
transform 1 0 52790 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_593
timestamp 1607639953
transform 1 0 55642 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_581
timestamp 1607639953
transform 1 0 54538 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_586
timestamp 1607639953
transform 1 0 54998 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_574
timestamp 1607639953
transform 1 0 53894 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1223
timestamp 1607639953
transform 1 0 54446 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_610
timestamp 1607639953
transform 1 0 57206 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_598
timestamp 1607639953
transform 1 0 56102 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_611
timestamp 1607639953
transform 1 0 57298 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_598
timestamp 1607639953
transform 1 0 56102 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1213
timestamp 1607639953
transform 1 0 57206 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _082_
timestamp 1607639953
transform 1 0 55826 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_100_622
timestamp 1607639953
transform 1 0 58310 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_623
timestamp 1607639953
transform 1 0 58402 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1607639953
transform -1 0 58862 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1607639953
transform -1 0 58862 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_15
timestamp 1607639953
transform 1 0 2466 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_3
timestamp 1607639953
transform 1 0 1362 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1607639953
transform 1 0 1086 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_44
timestamp 1607639953
transform 1 0 5134 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_32
timestamp 1607639953
transform 1 0 4030 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_27
timestamp 1607639953
transform 1 0 3570 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1224
timestamp 1607639953
transform 1 0 3938 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_63
timestamp 1607639953
transform 1 0 6882 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_56
timestamp 1607639953
transform 1 0 6238 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1225
timestamp 1607639953
transform 1 0 6790 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_87
timestamp 1607639953
transform 1 0 9090 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_75
timestamp 1607639953
transform 1 0 7986 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_106
timestamp 1607639953
transform 1 0 10838 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_94
timestamp 1607639953
transform 1 0 9734 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1226
timestamp 1607639953
transform 1 0 9642 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_125
timestamp 1607639953
transform 1 0 12586 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_118
timestamp 1607639953
transform 1 0 11942 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1227
timestamp 1607639953
transform 1 0 12494 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_149
timestamp 1607639953
transform 1 0 14794 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_137
timestamp 1607639953
transform 1 0 13690 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_168
timestamp 1607639953
transform 1 0 16542 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_156
timestamp 1607639953
transform 1 0 15438 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1228
timestamp 1607639953
transform 1 0 15346 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_187
timestamp 1607639953
transform 1 0 18290 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_180
timestamp 1607639953
transform 1 0 17646 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1229
timestamp 1607639953
transform 1 0 18198 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_218
timestamp 1607639953
transform 1 0 21142 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_211
timestamp 1607639953
transform 1 0 20498 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_199
timestamp 1607639953
transform 1 0 19394 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1230
timestamp 1607639953
transform 1 0 21050 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_242
timestamp 1607639953
transform 1 0 23350 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_230
timestamp 1607639953
transform 1 0 22246 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_261
timestamp 1607639953
transform 1 0 25098 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_249
timestamp 1607639953
transform 1 0 23994 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1231
timestamp 1607639953
transform 1 0 23902 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_280
timestamp 1607639953
transform 1 0 26846 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_273
timestamp 1607639953
transform 1 0 26202 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1232
timestamp 1607639953
transform 1 0 26754 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_304
timestamp 1607639953
transform 1 0 29054 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_292
timestamp 1607639953
transform 1 0 27950 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_323
timestamp 1607639953
transform 1 0 30802 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_311
timestamp 1607639953
transform 1 0 29698 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1233
timestamp 1607639953
transform 1 0 29606 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_342
timestamp 1607639953
transform 1 0 32550 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_335
timestamp 1607639953
transform 1 0 31906 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1234
timestamp 1607639953
transform 1 0 32458 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_373
timestamp 1607639953
transform 1 0 35402 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_366
timestamp 1607639953
transform 1 0 34758 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_354
timestamp 1607639953
transform 1 0 33654 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1235
timestamp 1607639953
transform 1 0 35310 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_385
timestamp 1607639953
transform 1 0 36506 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_416
timestamp 1607639953
transform 1 0 39358 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_404
timestamp 1607639953
transform 1 0 38254 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_397
timestamp 1607639953
transform 1 0 37610 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1236
timestamp 1607639953
transform 1 0 38162 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_435
timestamp 1607639953
transform 1 0 41106 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_428
timestamp 1607639953
transform 1 0 40462 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1237
timestamp 1607639953
transform 1 0 41014 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_459
timestamp 1607639953
transform 1 0 43314 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_447
timestamp 1607639953
transform 1 0 42210 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_478
timestamp 1607639953
transform 1 0 45062 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_466
timestamp 1607639953
transform 1 0 43958 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1238
timestamp 1607639953
transform 1 0 43866 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_497
timestamp 1607639953
transform 1 0 46810 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_490
timestamp 1607639953
transform 1 0 46166 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1239
timestamp 1607639953
transform 1 0 46718 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_528
timestamp 1607639953
transform 1 0 49662 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_521
timestamp 1607639953
transform 1 0 49018 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_509
timestamp 1607639953
transform 1 0 47914 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1240
timestamp 1607639953
transform 1 0 49570 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_540
timestamp 1607639953
transform 1 0 50766 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_571
timestamp 1607639953
transform 1 0 53618 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_559
timestamp 1607639953
transform 1 0 52514 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_552
timestamp 1607639953
transform 1 0 51870 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1241
timestamp 1607639953
transform 1 0 52422 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_590
timestamp 1607639953
transform 1 0 55366 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_583
timestamp 1607639953
transform 1 0 54722 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1242
timestamp 1607639953
transform 1 0 55274 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_614
timestamp 1607639953
transform 1 0 57574 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_602
timestamp 1607639953
transform 1 0 56470 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_621
timestamp 1607639953
transform 1 0 58218 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1243
timestamp 1607639953
transform 1 0 58126 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1607639953
transform -1 0 58862 0 1 57120
box -38 -48 314 592
<< labels >>
rlabel metal2 s 184 59200 240 60000 6 io_in[0]
port 0 nsew default input
rlabel metal2 s 15916 59200 15972 60000 6 io_in[10]
port 1 nsew default input
rlabel metal2 s 17480 59200 17536 60000 6 io_in[11]
port 2 nsew default input
rlabel metal2 s 19044 59200 19100 60000 6 io_in[12]
port 3 nsew default input
rlabel metal2 s 20700 59200 20756 60000 6 io_in[13]
port 4 nsew default input
rlabel metal2 s 22264 59200 22320 60000 6 io_in[14]
port 5 nsew default input
rlabel metal2 s 23828 59200 23884 60000 6 io_in[15]
port 6 nsew default input
rlabel metal2 s 25392 59200 25448 60000 6 io_in[16]
port 7 nsew default input
rlabel metal2 s 26956 59200 27012 60000 6 io_in[17]
port 8 nsew default input
rlabel metal2 s 28520 59200 28576 60000 6 io_in[18]
port 9 nsew default input
rlabel metal2 s 30176 59200 30232 60000 6 io_in[19]
port 10 nsew default input
rlabel metal2 s 1748 59200 1804 60000 6 io_in[1]
port 11 nsew default input
rlabel metal2 s 31740 59200 31796 60000 6 io_in[20]
port 12 nsew default input
rlabel metal2 s 33304 59200 33360 60000 6 io_in[21]
port 13 nsew default input
rlabel metal2 s 34868 59200 34924 60000 6 io_in[22]
port 14 nsew default input
rlabel metal2 s 36432 59200 36488 60000 6 io_in[23]
port 15 nsew default input
rlabel metal2 s 37996 59200 38052 60000 6 io_in[24]
port 16 nsew default input
rlabel metal2 s 39560 59200 39616 60000 6 io_in[25]
port 17 nsew default input
rlabel metal2 s 41216 59200 41272 60000 6 io_in[26]
port 18 nsew default input
rlabel metal2 s 42780 59200 42836 60000 6 io_in[27]
port 19 nsew default input
rlabel metal2 s 44344 59200 44400 60000 6 io_in[28]
port 20 nsew default input
rlabel metal2 s 45908 59200 45964 60000 6 io_in[29]
port 21 nsew default input
rlabel metal2 s 3312 59200 3368 60000 6 io_in[2]
port 22 nsew default input
rlabel metal2 s 47472 59200 47528 60000 6 io_in[30]
port 23 nsew default input
rlabel metal2 s 49036 59200 49092 60000 6 io_in[31]
port 24 nsew default input
rlabel metal2 s 50692 59200 50748 60000 6 io_in[32]
port 25 nsew default input
rlabel metal2 s 52256 59200 52312 60000 6 io_in[33]
port 26 nsew default input
rlabel metal2 s 53820 59200 53876 60000 6 io_in[34]
port 27 nsew default input
rlabel metal2 s 55384 59200 55440 60000 6 io_in[35]
port 28 nsew default input
rlabel metal2 s 56948 59200 57004 60000 6 io_in[36]
port 29 nsew default input
rlabel metal2 s 58512 59200 58568 60000 6 io_in[37]
port 30 nsew default input
rlabel metal2 s 4876 59200 4932 60000 6 io_in[3]
port 31 nsew default input
rlabel metal2 s 6440 59200 6496 60000 6 io_in[4]
port 32 nsew default input
rlabel metal2 s 8004 59200 8060 60000 6 io_in[5]
port 33 nsew default input
rlabel metal2 s 9568 59200 9624 60000 6 io_in[6]
port 34 nsew default input
rlabel metal2 s 11224 59200 11280 60000 6 io_in[7]
port 35 nsew default input
rlabel metal2 s 12788 59200 12844 60000 6 io_in[8]
port 36 nsew default input
rlabel metal2 s 14352 59200 14408 60000 6 io_in[9]
port 37 nsew default input
rlabel metal2 s 644 59200 700 60000 6 io_oeb[0]
port 38 nsew default tristate
rlabel metal2 s 16468 59200 16524 60000 6 io_oeb[10]
port 39 nsew default tristate
rlabel metal2 s 18032 59200 18088 60000 6 io_oeb[11]
port 40 nsew default tristate
rlabel metal2 s 19596 59200 19652 60000 6 io_oeb[12]
port 41 nsew default tristate
rlabel metal2 s 21160 59200 21216 60000 6 io_oeb[13]
port 42 nsew default tristate
rlabel metal2 s 22724 59200 22780 60000 6 io_oeb[14]
port 43 nsew default tristate
rlabel metal2 s 24380 59200 24436 60000 6 io_oeb[15]
port 44 nsew default tristate
rlabel metal2 s 25944 59200 26000 60000 6 io_oeb[16]
port 45 nsew default tristate
rlabel metal2 s 27508 59200 27564 60000 6 io_oeb[17]
port 46 nsew default tristate
rlabel metal2 s 29072 59200 29128 60000 6 io_oeb[18]
port 47 nsew default tristate
rlabel metal2 s 30636 59200 30692 60000 6 io_oeb[19]
port 48 nsew default tristate
rlabel metal2 s 2208 59200 2264 60000 6 io_oeb[1]
port 49 nsew default tristate
rlabel metal2 s 32200 59200 32256 60000 6 io_oeb[20]
port 50 nsew default tristate
rlabel metal2 s 33856 59200 33912 60000 6 io_oeb[21]
port 51 nsew default tristate
rlabel metal2 s 35420 59200 35476 60000 6 io_oeb[22]
port 52 nsew default tristate
rlabel metal2 s 36984 59200 37040 60000 6 io_oeb[23]
port 53 nsew default tristate
rlabel metal2 s 38548 59200 38604 60000 6 io_oeb[24]
port 54 nsew default tristate
rlabel metal2 s 40112 59200 40168 60000 6 io_oeb[25]
port 55 nsew default tristate
rlabel metal2 s 41676 59200 41732 60000 6 io_oeb[26]
port 56 nsew default tristate
rlabel metal2 s 43240 59200 43296 60000 6 io_oeb[27]
port 57 nsew default tristate
rlabel metal2 s 44896 59200 44952 60000 6 io_oeb[28]
port 58 nsew default tristate
rlabel metal2 s 46460 59200 46516 60000 6 io_oeb[29]
port 59 nsew default tristate
rlabel metal2 s 3864 59200 3920 60000 6 io_oeb[2]
port 60 nsew default tristate
rlabel metal2 s 48024 59200 48080 60000 6 io_oeb[30]
port 61 nsew default tristate
rlabel metal2 s 49588 59200 49644 60000 6 io_oeb[31]
port 62 nsew default tristate
rlabel metal2 s 51152 59200 51208 60000 6 io_oeb[32]
port 63 nsew default tristate
rlabel metal2 s 52716 59200 52772 60000 6 io_oeb[33]
port 64 nsew default tristate
rlabel metal2 s 54372 59200 54428 60000 6 io_oeb[34]
port 65 nsew default tristate
rlabel metal2 s 55936 59200 55992 60000 6 io_oeb[35]
port 66 nsew default tristate
rlabel metal2 s 57500 59200 57556 60000 6 io_oeb[36]
port 67 nsew default tristate
rlabel metal2 s 59064 59200 59120 60000 6 io_oeb[37]
port 68 nsew default tristate
rlabel metal2 s 5428 59200 5484 60000 6 io_oeb[3]
port 69 nsew default tristate
rlabel metal2 s 6992 59200 7048 60000 6 io_oeb[4]
port 70 nsew default tristate
rlabel metal2 s 8556 59200 8612 60000 6 io_oeb[5]
port 71 nsew default tristate
rlabel metal2 s 10120 59200 10176 60000 6 io_oeb[6]
port 72 nsew default tristate
rlabel metal2 s 11684 59200 11740 60000 6 io_oeb[7]
port 73 nsew default tristate
rlabel metal2 s 13248 59200 13304 60000 6 io_oeb[8]
port 74 nsew default tristate
rlabel metal2 s 14904 59200 14960 60000 6 io_oeb[9]
port 75 nsew default tristate
rlabel metal2 s 1196 59200 1252 60000 6 io_out[0]
port 76 nsew default tristate
rlabel metal2 s 17020 59200 17076 60000 6 io_out[10]
port 77 nsew default tristate
rlabel metal2 s 18584 59200 18640 60000 6 io_out[11]
port 78 nsew default tristate
rlabel metal2 s 20148 59200 20204 60000 6 io_out[12]
port 79 nsew default tristate
rlabel metal2 s 21712 59200 21768 60000 6 io_out[13]
port 80 nsew default tristate
rlabel metal2 s 23276 59200 23332 60000 6 io_out[14]
port 81 nsew default tristate
rlabel metal2 s 24840 59200 24896 60000 6 io_out[15]
port 82 nsew default tristate
rlabel metal2 s 26404 59200 26460 60000 6 io_out[16]
port 83 nsew default tristate
rlabel metal2 s 28060 59200 28116 60000 6 io_out[17]
port 84 nsew default tristate
rlabel metal2 s 29624 59200 29680 60000 6 io_out[18]
port 85 nsew default tristate
rlabel metal2 s 31188 59200 31244 60000 6 io_out[19]
port 86 nsew default tristate
rlabel metal2 s 2760 59200 2816 60000 6 io_out[1]
port 87 nsew default tristate
rlabel metal2 s 32752 59200 32808 60000 6 io_out[20]
port 88 nsew default tristate
rlabel metal2 s 34316 59200 34372 60000 6 io_out[21]
port 89 nsew default tristate
rlabel metal2 s 35880 59200 35936 60000 6 io_out[22]
port 90 nsew default tristate
rlabel metal2 s 37536 59200 37592 60000 6 io_out[23]
port 91 nsew default tristate
rlabel metal2 s 39100 59200 39156 60000 6 io_out[24]
port 92 nsew default tristate
rlabel metal2 s 40664 59200 40720 60000 6 io_out[25]
port 93 nsew default tristate
rlabel metal2 s 42228 59200 42284 60000 6 io_out[26]
port 94 nsew default tristate
rlabel metal2 s 43792 59200 43848 60000 6 io_out[27]
port 95 nsew default tristate
rlabel metal2 s 45356 59200 45412 60000 6 io_out[28]
port 96 nsew default tristate
rlabel metal2 s 47012 59200 47068 60000 6 io_out[29]
port 97 nsew default tristate
rlabel metal2 s 4324 59200 4380 60000 6 io_out[2]
port 98 nsew default tristate
rlabel metal2 s 48576 59200 48632 60000 6 io_out[30]
port 99 nsew default tristate
rlabel metal2 s 50140 59200 50196 60000 6 io_out[31]
port 100 nsew default tristate
rlabel metal2 s 51704 59200 51760 60000 6 io_out[32]
port 101 nsew default tristate
rlabel metal2 s 53268 59200 53324 60000 6 io_out[33]
port 102 nsew default tristate
rlabel metal2 s 54832 59200 54888 60000 6 io_out[34]
port 103 nsew default tristate
rlabel metal2 s 56396 59200 56452 60000 6 io_out[35]
port 104 nsew default tristate
rlabel metal2 s 58052 59200 58108 60000 6 io_out[36]
port 105 nsew default tristate
rlabel metal2 s 59616 59200 59672 60000 6 io_out[37]
port 106 nsew default tristate
rlabel metal2 s 5888 59200 5944 60000 6 io_out[3]
port 107 nsew default tristate
rlabel metal2 s 7544 59200 7600 60000 6 io_out[4]
port 108 nsew default tristate
rlabel metal2 s 9108 59200 9164 60000 6 io_out[5]
port 109 nsew default tristate
rlabel metal2 s 10672 59200 10728 60000 6 io_out[6]
port 110 nsew default tristate
rlabel metal2 s 12236 59200 12292 60000 6 io_out[7]
port 111 nsew default tristate
rlabel metal2 s 13800 59200 13856 60000 6 io_out[8]
port 112 nsew default tristate
rlabel metal2 s 15364 59200 15420 60000 6 io_out[9]
port 113 nsew default tristate
rlabel metal2 s 12972 0 13028 800 6 la_data_in[0]
port 114 nsew default input
rlabel metal2 s 49680 0 49736 800 6 la_data_in[100]
port 115 nsew default input
rlabel metal2 s 50048 0 50104 800 6 la_data_in[101]
port 116 nsew default input
rlabel metal2 s 50416 0 50472 800 6 la_data_in[102]
port 117 nsew default input
rlabel metal2 s 50784 0 50840 800 6 la_data_in[103]
port 118 nsew default input
rlabel metal2 s 51152 0 51208 800 6 la_data_in[104]
port 119 nsew default input
rlabel metal2 s 51520 0 51576 800 6 la_data_in[105]
port 120 nsew default input
rlabel metal2 s 51888 0 51944 800 6 la_data_in[106]
port 121 nsew default input
rlabel metal2 s 52256 0 52312 800 6 la_data_in[107]
port 122 nsew default input
rlabel metal2 s 52624 0 52680 800 6 la_data_in[108]
port 123 nsew default input
rlabel metal2 s 52992 0 53048 800 6 la_data_in[109]
port 124 nsew default input
rlabel metal2 s 16560 0 16616 800 6 la_data_in[10]
port 125 nsew default input
rlabel metal2 s 53360 0 53416 800 6 la_data_in[110]
port 126 nsew default input
rlabel metal2 s 53728 0 53784 800 6 la_data_in[111]
port 127 nsew default input
rlabel metal2 s 54096 0 54152 800 6 la_data_in[112]
port 128 nsew default input
rlabel metal2 s 54464 0 54520 800 6 la_data_in[113]
port 129 nsew default input
rlabel metal2 s 54832 0 54888 800 6 la_data_in[114]
port 130 nsew default input
rlabel metal2 s 55200 0 55256 800 6 la_data_in[115]
port 131 nsew default input
rlabel metal2 s 55568 0 55624 800 6 la_data_in[116]
port 132 nsew default input
rlabel metal2 s 55936 0 55992 800 6 la_data_in[117]
port 133 nsew default input
rlabel metal2 s 56304 0 56360 800 6 la_data_in[118]
port 134 nsew default input
rlabel metal2 s 56672 0 56728 800 6 la_data_in[119]
port 135 nsew default input
rlabel metal2 s 16928 0 16984 800 6 la_data_in[11]
port 136 nsew default input
rlabel metal2 s 57040 0 57096 800 6 la_data_in[120]
port 137 nsew default input
rlabel metal2 s 57408 0 57464 800 6 la_data_in[121]
port 138 nsew default input
rlabel metal2 s 57776 0 57832 800 6 la_data_in[122]
port 139 nsew default input
rlabel metal2 s 58144 0 58200 800 6 la_data_in[123]
port 140 nsew default input
rlabel metal2 s 58512 0 58568 800 6 la_data_in[124]
port 141 nsew default input
rlabel metal2 s 58880 0 58936 800 6 la_data_in[125]
port 142 nsew default input
rlabel metal2 s 59248 0 59304 800 6 la_data_in[126]
port 143 nsew default input
rlabel metal2 s 59616 0 59672 800 6 la_data_in[127]
port 144 nsew default input
rlabel metal2 s 17296 0 17352 800 6 la_data_in[12]
port 145 nsew default input
rlabel metal2 s 17664 0 17720 800 6 la_data_in[13]
port 146 nsew default input
rlabel metal2 s 18032 0 18088 800 6 la_data_in[14]
port 147 nsew default input
rlabel metal2 s 18400 0 18456 800 6 la_data_in[15]
port 148 nsew default input
rlabel metal2 s 18768 0 18824 800 6 la_data_in[16]
port 149 nsew default input
rlabel metal2 s 19136 0 19192 800 6 la_data_in[17]
port 150 nsew default input
rlabel metal2 s 19504 0 19560 800 6 la_data_in[18]
port 151 nsew default input
rlabel metal2 s 19872 0 19928 800 6 la_data_in[19]
port 152 nsew default input
rlabel metal2 s 13340 0 13396 800 6 la_data_in[1]
port 153 nsew default input
rlabel metal2 s 20240 0 20296 800 6 la_data_in[20]
port 154 nsew default input
rlabel metal2 s 20608 0 20664 800 6 la_data_in[21]
port 155 nsew default input
rlabel metal2 s 20976 0 21032 800 6 la_data_in[22]
port 156 nsew default input
rlabel metal2 s 21344 0 21400 800 6 la_data_in[23]
port 157 nsew default input
rlabel metal2 s 21712 0 21768 800 6 la_data_in[24]
port 158 nsew default input
rlabel metal2 s 22080 0 22136 800 6 la_data_in[25]
port 159 nsew default input
rlabel metal2 s 22448 0 22504 800 6 la_data_in[26]
port 160 nsew default input
rlabel metal2 s 22816 0 22872 800 6 la_data_in[27]
port 161 nsew default input
rlabel metal2 s 23184 0 23240 800 6 la_data_in[28]
port 162 nsew default input
rlabel metal2 s 23552 0 23608 800 6 la_data_in[29]
port 163 nsew default input
rlabel metal2 s 13708 0 13764 800 6 la_data_in[2]
port 164 nsew default input
rlabel metal2 s 23920 0 23976 800 6 la_data_in[30]
port 165 nsew default input
rlabel metal2 s 24288 0 24344 800 6 la_data_in[31]
port 166 nsew default input
rlabel metal2 s 24656 0 24712 800 6 la_data_in[32]
port 167 nsew default input
rlabel metal2 s 25024 0 25080 800 6 la_data_in[33]
port 168 nsew default input
rlabel metal2 s 25392 0 25448 800 6 la_data_in[34]
port 169 nsew default input
rlabel metal2 s 25760 0 25816 800 6 la_data_in[35]
port 170 nsew default input
rlabel metal2 s 26128 0 26184 800 6 la_data_in[36]
port 171 nsew default input
rlabel metal2 s 26496 0 26552 800 6 la_data_in[37]
port 172 nsew default input
rlabel metal2 s 26864 0 26920 800 6 la_data_in[38]
port 173 nsew default input
rlabel metal2 s 27232 0 27288 800 6 la_data_in[39]
port 174 nsew default input
rlabel metal2 s 14076 0 14132 800 6 la_data_in[3]
port 175 nsew default input
rlabel metal2 s 27600 0 27656 800 6 la_data_in[40]
port 176 nsew default input
rlabel metal2 s 27968 0 28024 800 6 la_data_in[41]
port 177 nsew default input
rlabel metal2 s 28336 0 28392 800 6 la_data_in[42]
port 178 nsew default input
rlabel metal2 s 28704 0 28760 800 6 la_data_in[43]
port 179 nsew default input
rlabel metal2 s 29072 0 29128 800 6 la_data_in[44]
port 180 nsew default input
rlabel metal2 s 29440 0 29496 800 6 la_data_in[45]
port 181 nsew default input
rlabel metal2 s 29808 0 29864 800 6 la_data_in[46]
port 182 nsew default input
rlabel metal2 s 30176 0 30232 800 6 la_data_in[47]
port 183 nsew default input
rlabel metal2 s 30544 0 30600 800 6 la_data_in[48]
port 184 nsew default input
rlabel metal2 s 30912 0 30968 800 6 la_data_in[49]
port 185 nsew default input
rlabel metal2 s 14444 0 14500 800 6 la_data_in[4]
port 186 nsew default input
rlabel metal2 s 31280 0 31336 800 6 la_data_in[50]
port 187 nsew default input
rlabel metal2 s 31648 0 31704 800 6 la_data_in[51]
port 188 nsew default input
rlabel metal2 s 32016 0 32072 800 6 la_data_in[52]
port 189 nsew default input
rlabel metal2 s 32384 0 32440 800 6 la_data_in[53]
port 190 nsew default input
rlabel metal2 s 32752 0 32808 800 6 la_data_in[54]
port 191 nsew default input
rlabel metal2 s 33120 0 33176 800 6 la_data_in[55]
port 192 nsew default input
rlabel metal2 s 33488 0 33544 800 6 la_data_in[56]
port 193 nsew default input
rlabel metal2 s 33856 0 33912 800 6 la_data_in[57]
port 194 nsew default input
rlabel metal2 s 34224 0 34280 800 6 la_data_in[58]
port 195 nsew default input
rlabel metal2 s 34592 0 34648 800 6 la_data_in[59]
port 196 nsew default input
rlabel metal2 s 14812 0 14868 800 6 la_data_in[5]
port 197 nsew default input
rlabel metal2 s 34960 0 35016 800 6 la_data_in[60]
port 198 nsew default input
rlabel metal2 s 35328 0 35384 800 6 la_data_in[61]
port 199 nsew default input
rlabel metal2 s 35696 0 35752 800 6 la_data_in[62]
port 200 nsew default input
rlabel metal2 s 36064 0 36120 800 6 la_data_in[63]
port 201 nsew default input
rlabel metal2 s 36432 0 36488 800 6 la_data_in[64]
port 202 nsew default input
rlabel metal2 s 36800 0 36856 800 6 la_data_in[65]
port 203 nsew default input
rlabel metal2 s 37168 0 37224 800 6 la_data_in[66]
port 204 nsew default input
rlabel metal2 s 37536 0 37592 800 6 la_data_in[67]
port 205 nsew default input
rlabel metal2 s 37904 0 37960 800 6 la_data_in[68]
port 206 nsew default input
rlabel metal2 s 38272 0 38328 800 6 la_data_in[69]
port 207 nsew default input
rlabel metal2 s 15088 0 15144 800 6 la_data_in[6]
port 208 nsew default input
rlabel metal2 s 38640 0 38696 800 6 la_data_in[70]
port 209 nsew default input
rlabel metal2 s 39008 0 39064 800 6 la_data_in[71]
port 210 nsew default input
rlabel metal2 s 39376 0 39432 800 6 la_data_in[72]
port 211 nsew default input
rlabel metal2 s 39744 0 39800 800 6 la_data_in[73]
port 212 nsew default input
rlabel metal2 s 40112 0 40168 800 6 la_data_in[74]
port 213 nsew default input
rlabel metal2 s 40480 0 40536 800 6 la_data_in[75]
port 214 nsew default input
rlabel metal2 s 40848 0 40904 800 6 la_data_in[76]
port 215 nsew default input
rlabel metal2 s 41216 0 41272 800 6 la_data_in[77]
port 216 nsew default input
rlabel metal2 s 41584 0 41640 800 6 la_data_in[78]
port 217 nsew default input
rlabel metal2 s 41952 0 42008 800 6 la_data_in[79]
port 218 nsew default input
rlabel metal2 s 15456 0 15512 800 6 la_data_in[7]
port 219 nsew default input
rlabel metal2 s 42320 0 42376 800 6 la_data_in[80]
port 220 nsew default input
rlabel metal2 s 42688 0 42744 800 6 la_data_in[81]
port 221 nsew default input
rlabel metal2 s 43056 0 43112 800 6 la_data_in[82]
port 222 nsew default input
rlabel metal2 s 43424 0 43480 800 6 la_data_in[83]
port 223 nsew default input
rlabel metal2 s 43792 0 43848 800 6 la_data_in[84]
port 224 nsew default input
rlabel metal2 s 44160 0 44216 800 6 la_data_in[85]
port 225 nsew default input
rlabel metal2 s 44528 0 44584 800 6 la_data_in[86]
port 226 nsew default input
rlabel metal2 s 44896 0 44952 800 6 la_data_in[87]
port 227 nsew default input
rlabel metal2 s 45264 0 45320 800 6 la_data_in[88]
port 228 nsew default input
rlabel metal2 s 45632 0 45688 800 6 la_data_in[89]
port 229 nsew default input
rlabel metal2 s 15824 0 15880 800 6 la_data_in[8]
port 230 nsew default input
rlabel metal2 s 46000 0 46056 800 6 la_data_in[90]
port 231 nsew default input
rlabel metal2 s 46368 0 46424 800 6 la_data_in[91]
port 232 nsew default input
rlabel metal2 s 46736 0 46792 800 6 la_data_in[92]
port 233 nsew default input
rlabel metal2 s 47104 0 47160 800 6 la_data_in[93]
port 234 nsew default input
rlabel metal2 s 47472 0 47528 800 6 la_data_in[94]
port 235 nsew default input
rlabel metal2 s 47840 0 47896 800 6 la_data_in[95]
port 236 nsew default input
rlabel metal2 s 48208 0 48264 800 6 la_data_in[96]
port 237 nsew default input
rlabel metal2 s 48576 0 48632 800 6 la_data_in[97]
port 238 nsew default input
rlabel metal2 s 48944 0 49000 800 6 la_data_in[98]
port 239 nsew default input
rlabel metal2 s 49312 0 49368 800 6 la_data_in[99]
port 240 nsew default input
rlabel metal2 s 16192 0 16248 800 6 la_data_in[9]
port 241 nsew default input
rlabel metal2 s 13064 0 13120 800 6 la_data_out[0]
port 242 nsew default tristate
rlabel metal2 s 49772 0 49828 800 6 la_data_out[100]
port 243 nsew default tristate
rlabel metal2 s 50140 0 50196 800 6 la_data_out[101]
port 244 nsew default tristate
rlabel metal2 s 50508 0 50564 800 6 la_data_out[102]
port 245 nsew default tristate
rlabel metal2 s 50876 0 50932 800 6 la_data_out[103]
port 246 nsew default tristate
rlabel metal2 s 51244 0 51300 800 6 la_data_out[104]
port 247 nsew default tristate
rlabel metal2 s 51612 0 51668 800 6 la_data_out[105]
port 248 nsew default tristate
rlabel metal2 s 51980 0 52036 800 6 la_data_out[106]
port 249 nsew default tristate
rlabel metal2 s 52348 0 52404 800 6 la_data_out[107]
port 250 nsew default tristate
rlabel metal2 s 52716 0 52772 800 6 la_data_out[108]
port 251 nsew default tristate
rlabel metal2 s 53084 0 53140 800 6 la_data_out[109]
port 252 nsew default tristate
rlabel metal2 s 16744 0 16800 800 6 la_data_out[10]
port 253 nsew default tristate
rlabel metal2 s 53452 0 53508 800 6 la_data_out[110]
port 254 nsew default tristate
rlabel metal2 s 53820 0 53876 800 6 la_data_out[111]
port 255 nsew default tristate
rlabel metal2 s 54188 0 54244 800 6 la_data_out[112]
port 256 nsew default tristate
rlabel metal2 s 54556 0 54612 800 6 la_data_out[113]
port 257 nsew default tristate
rlabel metal2 s 54924 0 54980 800 6 la_data_out[114]
port 258 nsew default tristate
rlabel metal2 s 55292 0 55348 800 6 la_data_out[115]
port 259 nsew default tristate
rlabel metal2 s 55660 0 55716 800 6 la_data_out[116]
port 260 nsew default tristate
rlabel metal2 s 56028 0 56084 800 6 la_data_out[117]
port 261 nsew default tristate
rlabel metal2 s 56396 0 56452 800 6 la_data_out[118]
port 262 nsew default tristate
rlabel metal2 s 56764 0 56820 800 6 la_data_out[119]
port 263 nsew default tristate
rlabel metal2 s 17112 0 17168 800 6 la_data_out[11]
port 264 nsew default tristate
rlabel metal2 s 57132 0 57188 800 6 la_data_out[120]
port 265 nsew default tristate
rlabel metal2 s 57500 0 57556 800 6 la_data_out[121]
port 266 nsew default tristate
rlabel metal2 s 57868 0 57924 800 6 la_data_out[122]
port 267 nsew default tristate
rlabel metal2 s 58236 0 58292 800 6 la_data_out[123]
port 268 nsew default tristate
rlabel metal2 s 58604 0 58660 800 6 la_data_out[124]
port 269 nsew default tristate
rlabel metal2 s 58972 0 59028 800 6 la_data_out[125]
port 270 nsew default tristate
rlabel metal2 s 59340 0 59396 800 6 la_data_out[126]
port 271 nsew default tristate
rlabel metal2 s 59708 0 59764 800 6 la_data_out[127]
port 272 nsew default tristate
rlabel metal2 s 17480 0 17536 800 6 la_data_out[12]
port 273 nsew default tristate
rlabel metal2 s 17848 0 17904 800 6 la_data_out[13]
port 274 nsew default tristate
rlabel metal2 s 18216 0 18272 800 6 la_data_out[14]
port 275 nsew default tristate
rlabel metal2 s 18584 0 18640 800 6 la_data_out[15]
port 276 nsew default tristate
rlabel metal2 s 18952 0 19008 800 6 la_data_out[16]
port 277 nsew default tristate
rlabel metal2 s 19320 0 19376 800 6 la_data_out[17]
port 278 nsew default tristate
rlabel metal2 s 19688 0 19744 800 6 la_data_out[18]
port 279 nsew default tristate
rlabel metal2 s 20056 0 20112 800 6 la_data_out[19]
port 280 nsew default tristate
rlabel metal2 s 13432 0 13488 800 6 la_data_out[1]
port 281 nsew default tristate
rlabel metal2 s 20424 0 20480 800 6 la_data_out[20]
port 282 nsew default tristate
rlabel metal2 s 20792 0 20848 800 6 la_data_out[21]
port 283 nsew default tristate
rlabel metal2 s 21160 0 21216 800 6 la_data_out[22]
port 284 nsew default tristate
rlabel metal2 s 21528 0 21584 800 6 la_data_out[23]
port 285 nsew default tristate
rlabel metal2 s 21896 0 21952 800 6 la_data_out[24]
port 286 nsew default tristate
rlabel metal2 s 22264 0 22320 800 6 la_data_out[25]
port 287 nsew default tristate
rlabel metal2 s 22632 0 22688 800 6 la_data_out[26]
port 288 nsew default tristate
rlabel metal2 s 23000 0 23056 800 6 la_data_out[27]
port 289 nsew default tristate
rlabel metal2 s 23368 0 23424 800 6 la_data_out[28]
port 290 nsew default tristate
rlabel metal2 s 23736 0 23792 800 6 la_data_out[29]
port 291 nsew default tristate
rlabel metal2 s 13800 0 13856 800 6 la_data_out[2]
port 292 nsew default tristate
rlabel metal2 s 24104 0 24160 800 6 la_data_out[30]
port 293 nsew default tristate
rlabel metal2 s 24472 0 24528 800 6 la_data_out[31]
port 294 nsew default tristate
rlabel metal2 s 24840 0 24896 800 6 la_data_out[32]
port 295 nsew default tristate
rlabel metal2 s 25208 0 25264 800 6 la_data_out[33]
port 296 nsew default tristate
rlabel metal2 s 25576 0 25632 800 6 la_data_out[34]
port 297 nsew default tristate
rlabel metal2 s 25944 0 26000 800 6 la_data_out[35]
port 298 nsew default tristate
rlabel metal2 s 26312 0 26368 800 6 la_data_out[36]
port 299 nsew default tristate
rlabel metal2 s 26680 0 26736 800 6 la_data_out[37]
port 300 nsew default tristate
rlabel metal2 s 27048 0 27104 800 6 la_data_out[38]
port 301 nsew default tristate
rlabel metal2 s 27416 0 27472 800 6 la_data_out[39]
port 302 nsew default tristate
rlabel metal2 s 14168 0 14224 800 6 la_data_out[3]
port 303 nsew default tristate
rlabel metal2 s 27784 0 27840 800 6 la_data_out[40]
port 304 nsew default tristate
rlabel metal2 s 28152 0 28208 800 6 la_data_out[41]
port 305 nsew default tristate
rlabel metal2 s 28520 0 28576 800 6 la_data_out[42]
port 306 nsew default tristate
rlabel metal2 s 28888 0 28944 800 6 la_data_out[43]
port 307 nsew default tristate
rlabel metal2 s 29256 0 29312 800 6 la_data_out[44]
port 308 nsew default tristate
rlabel metal2 s 29624 0 29680 800 6 la_data_out[45]
port 309 nsew default tristate
rlabel metal2 s 29992 0 30048 800 6 la_data_out[46]
port 310 nsew default tristate
rlabel metal2 s 30268 0 30324 800 6 la_data_out[47]
port 311 nsew default tristate
rlabel metal2 s 30636 0 30692 800 6 la_data_out[48]
port 312 nsew default tristate
rlabel metal2 s 31004 0 31060 800 6 la_data_out[49]
port 313 nsew default tristate
rlabel metal2 s 14536 0 14592 800 6 la_data_out[4]
port 314 nsew default tristate
rlabel metal2 s 31372 0 31428 800 6 la_data_out[50]
port 315 nsew default tristate
rlabel metal2 s 31740 0 31796 800 6 la_data_out[51]
port 316 nsew default tristate
rlabel metal2 s 32108 0 32164 800 6 la_data_out[52]
port 317 nsew default tristate
rlabel metal2 s 32476 0 32532 800 6 la_data_out[53]
port 318 nsew default tristate
rlabel metal2 s 32844 0 32900 800 6 la_data_out[54]
port 319 nsew default tristate
rlabel metal2 s 33212 0 33268 800 6 la_data_out[55]
port 320 nsew default tristate
rlabel metal2 s 33580 0 33636 800 6 la_data_out[56]
port 321 nsew default tristate
rlabel metal2 s 33948 0 34004 800 6 la_data_out[57]
port 322 nsew default tristate
rlabel metal2 s 34316 0 34372 800 6 la_data_out[58]
port 323 nsew default tristate
rlabel metal2 s 34684 0 34740 800 6 la_data_out[59]
port 324 nsew default tristate
rlabel metal2 s 14904 0 14960 800 6 la_data_out[5]
port 325 nsew default tristate
rlabel metal2 s 35052 0 35108 800 6 la_data_out[60]
port 326 nsew default tristate
rlabel metal2 s 35420 0 35476 800 6 la_data_out[61]
port 327 nsew default tristate
rlabel metal2 s 35788 0 35844 800 6 la_data_out[62]
port 328 nsew default tristate
rlabel metal2 s 36156 0 36212 800 6 la_data_out[63]
port 329 nsew default tristate
rlabel metal2 s 36524 0 36580 800 6 la_data_out[64]
port 330 nsew default tristate
rlabel metal2 s 36892 0 36948 800 6 la_data_out[65]
port 331 nsew default tristate
rlabel metal2 s 37260 0 37316 800 6 la_data_out[66]
port 332 nsew default tristate
rlabel metal2 s 37628 0 37684 800 6 la_data_out[67]
port 333 nsew default tristate
rlabel metal2 s 37996 0 38052 800 6 la_data_out[68]
port 334 nsew default tristate
rlabel metal2 s 38364 0 38420 800 6 la_data_out[69]
port 335 nsew default tristate
rlabel metal2 s 15272 0 15328 800 6 la_data_out[6]
port 336 nsew default tristate
rlabel metal2 s 38732 0 38788 800 6 la_data_out[70]
port 337 nsew default tristate
rlabel metal2 s 39100 0 39156 800 6 la_data_out[71]
port 338 nsew default tristate
rlabel metal2 s 39468 0 39524 800 6 la_data_out[72]
port 339 nsew default tristate
rlabel metal2 s 39836 0 39892 800 6 la_data_out[73]
port 340 nsew default tristate
rlabel metal2 s 40204 0 40260 800 6 la_data_out[74]
port 341 nsew default tristate
rlabel metal2 s 40572 0 40628 800 6 la_data_out[75]
port 342 nsew default tristate
rlabel metal2 s 40940 0 40996 800 6 la_data_out[76]
port 343 nsew default tristate
rlabel metal2 s 41308 0 41364 800 6 la_data_out[77]
port 344 nsew default tristate
rlabel metal2 s 41676 0 41732 800 6 la_data_out[78]
port 345 nsew default tristate
rlabel metal2 s 42044 0 42100 800 6 la_data_out[79]
port 346 nsew default tristate
rlabel metal2 s 15640 0 15696 800 6 la_data_out[7]
port 347 nsew default tristate
rlabel metal2 s 42412 0 42468 800 6 la_data_out[80]
port 348 nsew default tristate
rlabel metal2 s 42780 0 42836 800 6 la_data_out[81]
port 349 nsew default tristate
rlabel metal2 s 43148 0 43204 800 6 la_data_out[82]
port 350 nsew default tristate
rlabel metal2 s 43516 0 43572 800 6 la_data_out[83]
port 351 nsew default tristate
rlabel metal2 s 43884 0 43940 800 6 la_data_out[84]
port 352 nsew default tristate
rlabel metal2 s 44252 0 44308 800 6 la_data_out[85]
port 353 nsew default tristate
rlabel metal2 s 44620 0 44676 800 6 la_data_out[86]
port 354 nsew default tristate
rlabel metal2 s 44988 0 45044 800 6 la_data_out[87]
port 355 nsew default tristate
rlabel metal2 s 45356 0 45412 800 6 la_data_out[88]
port 356 nsew default tristate
rlabel metal2 s 45724 0 45780 800 6 la_data_out[89]
port 357 nsew default tristate
rlabel metal2 s 16008 0 16064 800 6 la_data_out[8]
port 358 nsew default tristate
rlabel metal2 s 46092 0 46148 800 6 la_data_out[90]
port 359 nsew default tristate
rlabel metal2 s 46460 0 46516 800 6 la_data_out[91]
port 360 nsew default tristate
rlabel metal2 s 46828 0 46884 800 6 la_data_out[92]
port 361 nsew default tristate
rlabel metal2 s 47196 0 47252 800 6 la_data_out[93]
port 362 nsew default tristate
rlabel metal2 s 47564 0 47620 800 6 la_data_out[94]
port 363 nsew default tristate
rlabel metal2 s 47932 0 47988 800 6 la_data_out[95]
port 364 nsew default tristate
rlabel metal2 s 48300 0 48356 800 6 la_data_out[96]
port 365 nsew default tristate
rlabel metal2 s 48668 0 48724 800 6 la_data_out[97]
port 366 nsew default tristate
rlabel metal2 s 49036 0 49092 800 6 la_data_out[98]
port 367 nsew default tristate
rlabel metal2 s 49404 0 49460 800 6 la_data_out[99]
port 368 nsew default tristate
rlabel metal2 s 16376 0 16432 800 6 la_data_out[9]
port 369 nsew default tristate
rlabel metal2 s 13156 0 13212 800 6 la_oen[0]
port 370 nsew default input
rlabel metal2 s 49864 0 49920 800 6 la_oen[100]
port 371 nsew default input
rlabel metal2 s 50232 0 50288 800 6 la_oen[101]
port 372 nsew default input
rlabel metal2 s 50600 0 50656 800 6 la_oen[102]
port 373 nsew default input
rlabel metal2 s 50968 0 51024 800 6 la_oen[103]
port 374 nsew default input
rlabel metal2 s 51336 0 51392 800 6 la_oen[104]
port 375 nsew default input
rlabel metal2 s 51704 0 51760 800 6 la_oen[105]
port 376 nsew default input
rlabel metal2 s 52072 0 52128 800 6 la_oen[106]
port 377 nsew default input
rlabel metal2 s 52440 0 52496 800 6 la_oen[107]
port 378 nsew default input
rlabel metal2 s 52808 0 52864 800 6 la_oen[108]
port 379 nsew default input
rlabel metal2 s 53176 0 53232 800 6 la_oen[109]
port 380 nsew default input
rlabel metal2 s 16836 0 16892 800 6 la_oen[10]
port 381 nsew default input
rlabel metal2 s 53544 0 53600 800 6 la_oen[110]
port 382 nsew default input
rlabel metal2 s 53912 0 53968 800 6 la_oen[111]
port 383 nsew default input
rlabel metal2 s 54280 0 54336 800 6 la_oen[112]
port 384 nsew default input
rlabel metal2 s 54648 0 54704 800 6 la_oen[113]
port 385 nsew default input
rlabel metal2 s 55016 0 55072 800 6 la_oen[114]
port 386 nsew default input
rlabel metal2 s 55384 0 55440 800 6 la_oen[115]
port 387 nsew default input
rlabel metal2 s 55752 0 55808 800 6 la_oen[116]
port 388 nsew default input
rlabel metal2 s 56120 0 56176 800 6 la_oen[117]
port 389 nsew default input
rlabel metal2 s 56488 0 56544 800 6 la_oen[118]
port 390 nsew default input
rlabel metal2 s 56856 0 56912 800 6 la_oen[119]
port 391 nsew default input
rlabel metal2 s 17204 0 17260 800 6 la_oen[11]
port 392 nsew default input
rlabel metal2 s 57224 0 57280 800 6 la_oen[120]
port 393 nsew default input
rlabel metal2 s 57592 0 57648 800 6 la_oen[121]
port 394 nsew default input
rlabel metal2 s 57960 0 58016 800 6 la_oen[122]
port 395 nsew default input
rlabel metal2 s 58328 0 58384 800 6 la_oen[123]
port 396 nsew default input
rlabel metal2 s 58696 0 58752 800 6 la_oen[124]
port 397 nsew default input
rlabel metal2 s 59064 0 59120 800 6 la_oen[125]
port 398 nsew default input
rlabel metal2 s 59432 0 59488 800 6 la_oen[126]
port 399 nsew default input
rlabel metal2 s 59800 0 59856 800 6 la_oen[127]
port 400 nsew default input
rlabel metal2 s 17572 0 17628 800 6 la_oen[12]
port 401 nsew default input
rlabel metal2 s 17940 0 17996 800 6 la_oen[13]
port 402 nsew default input
rlabel metal2 s 18308 0 18364 800 6 la_oen[14]
port 403 nsew default input
rlabel metal2 s 18676 0 18732 800 6 la_oen[15]
port 404 nsew default input
rlabel metal2 s 19044 0 19100 800 6 la_oen[16]
port 405 nsew default input
rlabel metal2 s 19412 0 19468 800 6 la_oen[17]
port 406 nsew default input
rlabel metal2 s 19780 0 19836 800 6 la_oen[18]
port 407 nsew default input
rlabel metal2 s 20148 0 20204 800 6 la_oen[19]
port 408 nsew default input
rlabel metal2 s 13524 0 13580 800 6 la_oen[1]
port 409 nsew default input
rlabel metal2 s 20516 0 20572 800 6 la_oen[20]
port 410 nsew default input
rlabel metal2 s 20884 0 20940 800 6 la_oen[21]
port 411 nsew default input
rlabel metal2 s 21252 0 21308 800 6 la_oen[22]
port 412 nsew default input
rlabel metal2 s 21620 0 21676 800 6 la_oen[23]
port 413 nsew default input
rlabel metal2 s 21988 0 22044 800 6 la_oen[24]
port 414 nsew default input
rlabel metal2 s 22356 0 22412 800 6 la_oen[25]
port 415 nsew default input
rlabel metal2 s 22724 0 22780 800 6 la_oen[26]
port 416 nsew default input
rlabel metal2 s 23092 0 23148 800 6 la_oen[27]
port 417 nsew default input
rlabel metal2 s 23460 0 23516 800 6 la_oen[28]
port 418 nsew default input
rlabel metal2 s 23828 0 23884 800 6 la_oen[29]
port 419 nsew default input
rlabel metal2 s 13892 0 13948 800 6 la_oen[2]
port 420 nsew default input
rlabel metal2 s 24196 0 24252 800 6 la_oen[30]
port 421 nsew default input
rlabel metal2 s 24564 0 24620 800 6 la_oen[31]
port 422 nsew default input
rlabel metal2 s 24932 0 24988 800 6 la_oen[32]
port 423 nsew default input
rlabel metal2 s 25300 0 25356 800 6 la_oen[33]
port 424 nsew default input
rlabel metal2 s 25668 0 25724 800 6 la_oen[34]
port 425 nsew default input
rlabel metal2 s 26036 0 26092 800 6 la_oen[35]
port 426 nsew default input
rlabel metal2 s 26404 0 26460 800 6 la_oen[36]
port 427 nsew default input
rlabel metal2 s 26772 0 26828 800 6 la_oen[37]
port 428 nsew default input
rlabel metal2 s 27140 0 27196 800 6 la_oen[38]
port 429 nsew default input
rlabel metal2 s 27508 0 27564 800 6 la_oen[39]
port 430 nsew default input
rlabel metal2 s 14260 0 14316 800 6 la_oen[3]
port 431 nsew default input
rlabel metal2 s 27876 0 27932 800 6 la_oen[40]
port 432 nsew default input
rlabel metal2 s 28244 0 28300 800 6 la_oen[41]
port 433 nsew default input
rlabel metal2 s 28612 0 28668 800 6 la_oen[42]
port 434 nsew default input
rlabel metal2 s 28980 0 29036 800 6 la_oen[43]
port 435 nsew default input
rlabel metal2 s 29348 0 29404 800 6 la_oen[44]
port 436 nsew default input
rlabel metal2 s 29716 0 29772 800 6 la_oen[45]
port 437 nsew default input
rlabel metal2 s 30084 0 30140 800 6 la_oen[46]
port 438 nsew default input
rlabel metal2 s 30452 0 30508 800 6 la_oen[47]
port 439 nsew default input
rlabel metal2 s 30820 0 30876 800 6 la_oen[48]
port 440 nsew default input
rlabel metal2 s 31188 0 31244 800 6 la_oen[49]
port 441 nsew default input
rlabel metal2 s 14628 0 14684 800 6 la_oen[4]
port 442 nsew default input
rlabel metal2 s 31556 0 31612 800 6 la_oen[50]
port 443 nsew default input
rlabel metal2 s 31924 0 31980 800 6 la_oen[51]
port 444 nsew default input
rlabel metal2 s 32292 0 32348 800 6 la_oen[52]
port 445 nsew default input
rlabel metal2 s 32660 0 32716 800 6 la_oen[53]
port 446 nsew default input
rlabel metal2 s 33028 0 33084 800 6 la_oen[54]
port 447 nsew default input
rlabel metal2 s 33396 0 33452 800 6 la_oen[55]
port 448 nsew default input
rlabel metal2 s 33764 0 33820 800 6 la_oen[56]
port 449 nsew default input
rlabel metal2 s 34132 0 34188 800 6 la_oen[57]
port 450 nsew default input
rlabel metal2 s 34500 0 34556 800 6 la_oen[58]
port 451 nsew default input
rlabel metal2 s 34868 0 34924 800 6 la_oen[59]
port 452 nsew default input
rlabel metal2 s 14996 0 15052 800 6 la_oen[5]
port 453 nsew default input
rlabel metal2 s 35236 0 35292 800 6 la_oen[60]
port 454 nsew default input
rlabel metal2 s 35604 0 35660 800 6 la_oen[61]
port 455 nsew default input
rlabel metal2 s 35972 0 36028 800 6 la_oen[62]
port 456 nsew default input
rlabel metal2 s 36340 0 36396 800 6 la_oen[63]
port 457 nsew default input
rlabel metal2 s 36708 0 36764 800 6 la_oen[64]
port 458 nsew default input
rlabel metal2 s 37076 0 37132 800 6 la_oen[65]
port 459 nsew default input
rlabel metal2 s 37444 0 37500 800 6 la_oen[66]
port 460 nsew default input
rlabel metal2 s 37812 0 37868 800 6 la_oen[67]
port 461 nsew default input
rlabel metal2 s 38180 0 38236 800 6 la_oen[68]
port 462 nsew default input
rlabel metal2 s 38548 0 38604 800 6 la_oen[69]
port 463 nsew default input
rlabel metal2 s 15364 0 15420 800 6 la_oen[6]
port 464 nsew default input
rlabel metal2 s 38916 0 38972 800 6 la_oen[70]
port 465 nsew default input
rlabel metal2 s 39284 0 39340 800 6 la_oen[71]
port 466 nsew default input
rlabel metal2 s 39652 0 39708 800 6 la_oen[72]
port 467 nsew default input
rlabel metal2 s 40020 0 40076 800 6 la_oen[73]
port 468 nsew default input
rlabel metal2 s 40388 0 40444 800 6 la_oen[74]
port 469 nsew default input
rlabel metal2 s 40756 0 40812 800 6 la_oen[75]
port 470 nsew default input
rlabel metal2 s 41124 0 41180 800 6 la_oen[76]
port 471 nsew default input
rlabel metal2 s 41492 0 41548 800 6 la_oen[77]
port 472 nsew default input
rlabel metal2 s 41860 0 41916 800 6 la_oen[78]
port 473 nsew default input
rlabel metal2 s 42228 0 42284 800 6 la_oen[79]
port 474 nsew default input
rlabel metal2 s 15732 0 15788 800 6 la_oen[7]
port 475 nsew default input
rlabel metal2 s 42596 0 42652 800 6 la_oen[80]
port 476 nsew default input
rlabel metal2 s 42964 0 43020 800 6 la_oen[81]
port 477 nsew default input
rlabel metal2 s 43332 0 43388 800 6 la_oen[82]
port 478 nsew default input
rlabel metal2 s 43700 0 43756 800 6 la_oen[83]
port 479 nsew default input
rlabel metal2 s 44068 0 44124 800 6 la_oen[84]
port 480 nsew default input
rlabel metal2 s 44436 0 44492 800 6 la_oen[85]
port 481 nsew default input
rlabel metal2 s 44804 0 44860 800 6 la_oen[86]
port 482 nsew default input
rlabel metal2 s 45080 0 45136 800 6 la_oen[87]
port 483 nsew default input
rlabel metal2 s 45448 0 45504 800 6 la_oen[88]
port 484 nsew default input
rlabel metal2 s 45816 0 45872 800 6 la_oen[89]
port 485 nsew default input
rlabel metal2 s 16100 0 16156 800 6 la_oen[8]
port 486 nsew default input
rlabel metal2 s 46184 0 46240 800 6 la_oen[90]
port 487 nsew default input
rlabel metal2 s 46552 0 46608 800 6 la_oen[91]
port 488 nsew default input
rlabel metal2 s 46920 0 46976 800 6 la_oen[92]
port 489 nsew default input
rlabel metal2 s 47288 0 47344 800 6 la_oen[93]
port 490 nsew default input
rlabel metal2 s 47656 0 47712 800 6 la_oen[94]
port 491 nsew default input
rlabel metal2 s 48024 0 48080 800 6 la_oen[95]
port 492 nsew default input
rlabel metal2 s 48392 0 48448 800 6 la_oen[96]
port 493 nsew default input
rlabel metal2 s 48760 0 48816 800 6 la_oen[97]
port 494 nsew default input
rlabel metal2 s 49128 0 49184 800 6 la_oen[98]
port 495 nsew default input
rlabel metal2 s 49496 0 49552 800 6 la_oen[99]
port 496 nsew default input
rlabel metal2 s 16468 0 16524 800 6 la_oen[9]
port 497 nsew default input
rlabel metal2 s 0 0 56 800 6 wb_clk_i
port 498 nsew default input
rlabel metal2 s 92 0 148 800 6 wb_rst_i
port 499 nsew default input
rlabel metal2 s 184 0 240 800 6 wbs_ack_o
port 500 nsew default tristate
rlabel metal2 s 644 0 700 800 6 wbs_adr_i[0]
port 501 nsew default input
rlabel metal2 s 4876 0 4932 800 6 wbs_adr_i[10]
port 502 nsew default input
rlabel metal2 s 5244 0 5300 800 6 wbs_adr_i[11]
port 503 nsew default input
rlabel metal2 s 5612 0 5668 800 6 wbs_adr_i[12]
port 504 nsew default input
rlabel metal2 s 5980 0 6036 800 6 wbs_adr_i[13]
port 505 nsew default input
rlabel metal2 s 6348 0 6404 800 6 wbs_adr_i[14]
port 506 nsew default input
rlabel metal2 s 6716 0 6772 800 6 wbs_adr_i[15]
port 507 nsew default input
rlabel metal2 s 7084 0 7140 800 6 wbs_adr_i[16]
port 508 nsew default input
rlabel metal2 s 7452 0 7508 800 6 wbs_adr_i[17]
port 509 nsew default input
rlabel metal2 s 7820 0 7876 800 6 wbs_adr_i[18]
port 510 nsew default input
rlabel metal2 s 8188 0 8244 800 6 wbs_adr_i[19]
port 511 nsew default input
rlabel metal2 s 1196 0 1252 800 6 wbs_adr_i[1]
port 512 nsew default input
rlabel metal2 s 8556 0 8612 800 6 wbs_adr_i[20]
port 513 nsew default input
rlabel metal2 s 8924 0 8980 800 6 wbs_adr_i[21]
port 514 nsew default input
rlabel metal2 s 9292 0 9348 800 6 wbs_adr_i[22]
port 515 nsew default input
rlabel metal2 s 9660 0 9716 800 6 wbs_adr_i[23]
port 516 nsew default input
rlabel metal2 s 10028 0 10084 800 6 wbs_adr_i[24]
port 517 nsew default input
rlabel metal2 s 10396 0 10452 800 6 wbs_adr_i[25]
port 518 nsew default input
rlabel metal2 s 10764 0 10820 800 6 wbs_adr_i[26]
port 519 nsew default input
rlabel metal2 s 11132 0 11188 800 6 wbs_adr_i[27]
port 520 nsew default input
rlabel metal2 s 11500 0 11556 800 6 wbs_adr_i[28]
port 521 nsew default input
rlabel metal2 s 11868 0 11924 800 6 wbs_adr_i[29]
port 522 nsew default input
rlabel metal2 s 1656 0 1712 800 6 wbs_adr_i[2]
port 523 nsew default input
rlabel metal2 s 12236 0 12292 800 6 wbs_adr_i[30]
port 524 nsew default input
rlabel metal2 s 12604 0 12660 800 6 wbs_adr_i[31]
port 525 nsew default input
rlabel metal2 s 2116 0 2172 800 6 wbs_adr_i[3]
port 526 nsew default input
rlabel metal2 s 2668 0 2724 800 6 wbs_adr_i[4]
port 527 nsew default input
rlabel metal2 s 3036 0 3092 800 6 wbs_adr_i[5]
port 528 nsew default input
rlabel metal2 s 3404 0 3460 800 6 wbs_adr_i[6]
port 529 nsew default input
rlabel metal2 s 3772 0 3828 800 6 wbs_adr_i[7]
port 530 nsew default input
rlabel metal2 s 4140 0 4196 800 6 wbs_adr_i[8]
port 531 nsew default input
rlabel metal2 s 4508 0 4564 800 6 wbs_adr_i[9]
port 532 nsew default input
rlabel metal2 s 276 0 332 800 6 wbs_cyc_i
port 533 nsew default input
rlabel metal2 s 828 0 884 800 6 wbs_dat_i[0]
port 534 nsew default input
rlabel metal2 s 4968 0 5024 800 6 wbs_dat_i[10]
port 535 nsew default input
rlabel metal2 s 5336 0 5392 800 6 wbs_dat_i[11]
port 536 nsew default input
rlabel metal2 s 5704 0 5760 800 6 wbs_dat_i[12]
port 537 nsew default input
rlabel metal2 s 6072 0 6128 800 6 wbs_dat_i[13]
port 538 nsew default input
rlabel metal2 s 6440 0 6496 800 6 wbs_dat_i[14]
port 539 nsew default input
rlabel metal2 s 6808 0 6864 800 6 wbs_dat_i[15]
port 540 nsew default input
rlabel metal2 s 7176 0 7232 800 6 wbs_dat_i[16]
port 541 nsew default input
rlabel metal2 s 7544 0 7600 800 6 wbs_dat_i[17]
port 542 nsew default input
rlabel metal2 s 7912 0 7968 800 6 wbs_dat_i[18]
port 543 nsew default input
rlabel metal2 s 8280 0 8336 800 6 wbs_dat_i[19]
port 544 nsew default input
rlabel metal2 s 1288 0 1344 800 6 wbs_dat_i[1]
port 545 nsew default input
rlabel metal2 s 8648 0 8704 800 6 wbs_dat_i[20]
port 546 nsew default input
rlabel metal2 s 9016 0 9072 800 6 wbs_dat_i[21]
port 547 nsew default input
rlabel metal2 s 9384 0 9440 800 6 wbs_dat_i[22]
port 548 nsew default input
rlabel metal2 s 9752 0 9808 800 6 wbs_dat_i[23]
port 549 nsew default input
rlabel metal2 s 10120 0 10176 800 6 wbs_dat_i[24]
port 550 nsew default input
rlabel metal2 s 10488 0 10544 800 6 wbs_dat_i[25]
port 551 nsew default input
rlabel metal2 s 10856 0 10912 800 6 wbs_dat_i[26]
port 552 nsew default input
rlabel metal2 s 11224 0 11280 800 6 wbs_dat_i[27]
port 553 nsew default input
rlabel metal2 s 11592 0 11648 800 6 wbs_dat_i[28]
port 554 nsew default input
rlabel metal2 s 11960 0 12016 800 6 wbs_dat_i[29]
port 555 nsew default input
rlabel metal2 s 1748 0 1804 800 6 wbs_dat_i[2]
port 556 nsew default input
rlabel metal2 s 12328 0 12384 800 6 wbs_dat_i[30]
port 557 nsew default input
rlabel metal2 s 12696 0 12752 800 6 wbs_dat_i[31]
port 558 nsew default input
rlabel metal2 s 2300 0 2356 800 6 wbs_dat_i[3]
port 559 nsew default input
rlabel metal2 s 2760 0 2816 800 6 wbs_dat_i[4]
port 560 nsew default input
rlabel metal2 s 3128 0 3184 800 6 wbs_dat_i[5]
port 561 nsew default input
rlabel metal2 s 3496 0 3552 800 6 wbs_dat_i[6]
port 562 nsew default input
rlabel metal2 s 3864 0 3920 800 6 wbs_dat_i[7]
port 563 nsew default input
rlabel metal2 s 4232 0 4288 800 6 wbs_dat_i[8]
port 564 nsew default input
rlabel metal2 s 4600 0 4656 800 6 wbs_dat_i[9]
port 565 nsew default input
rlabel metal2 s 920 0 976 800 6 wbs_dat_o[0]
port 566 nsew default tristate
rlabel metal2 s 5060 0 5116 800 6 wbs_dat_o[10]
port 567 nsew default tristate
rlabel metal2 s 5428 0 5484 800 6 wbs_dat_o[11]
port 568 nsew default tristate
rlabel metal2 s 5796 0 5852 800 6 wbs_dat_o[12]
port 569 nsew default tristate
rlabel metal2 s 6164 0 6220 800 6 wbs_dat_o[13]
port 570 nsew default tristate
rlabel metal2 s 6532 0 6588 800 6 wbs_dat_o[14]
port 571 nsew default tristate
rlabel metal2 s 6900 0 6956 800 6 wbs_dat_o[15]
port 572 nsew default tristate
rlabel metal2 s 7268 0 7324 800 6 wbs_dat_o[16]
port 573 nsew default tristate
rlabel metal2 s 7636 0 7692 800 6 wbs_dat_o[17]
port 574 nsew default tristate
rlabel metal2 s 8004 0 8060 800 6 wbs_dat_o[18]
port 575 nsew default tristate
rlabel metal2 s 8372 0 8428 800 6 wbs_dat_o[19]
port 576 nsew default tristate
rlabel metal2 s 1380 0 1436 800 6 wbs_dat_o[1]
port 577 nsew default tristate
rlabel metal2 s 8740 0 8796 800 6 wbs_dat_o[20]
port 578 nsew default tristate
rlabel metal2 s 9108 0 9164 800 6 wbs_dat_o[21]
port 579 nsew default tristate
rlabel metal2 s 9476 0 9532 800 6 wbs_dat_o[22]
port 580 nsew default tristate
rlabel metal2 s 9844 0 9900 800 6 wbs_dat_o[23]
port 581 nsew default tristate
rlabel metal2 s 10212 0 10268 800 6 wbs_dat_o[24]
port 582 nsew default tristate
rlabel metal2 s 10580 0 10636 800 6 wbs_dat_o[25]
port 583 nsew default tristate
rlabel metal2 s 10948 0 11004 800 6 wbs_dat_o[26]
port 584 nsew default tristate
rlabel metal2 s 11316 0 11372 800 6 wbs_dat_o[27]
port 585 nsew default tristate
rlabel metal2 s 11684 0 11740 800 6 wbs_dat_o[28]
port 586 nsew default tristate
rlabel metal2 s 12052 0 12108 800 6 wbs_dat_o[29]
port 587 nsew default tristate
rlabel metal2 s 1932 0 1988 800 6 wbs_dat_o[2]
port 588 nsew default tristate
rlabel metal2 s 12420 0 12476 800 6 wbs_dat_o[30]
port 589 nsew default tristate
rlabel metal2 s 12788 0 12844 800 6 wbs_dat_o[31]
port 590 nsew default tristate
rlabel metal2 s 2392 0 2448 800 6 wbs_dat_o[3]
port 591 nsew default tristate
rlabel metal2 s 2852 0 2908 800 6 wbs_dat_o[4]
port 592 nsew default tristate
rlabel metal2 s 3220 0 3276 800 6 wbs_dat_o[5]
port 593 nsew default tristate
rlabel metal2 s 3588 0 3644 800 6 wbs_dat_o[6]
port 594 nsew default tristate
rlabel metal2 s 3956 0 4012 800 6 wbs_dat_o[7]
port 595 nsew default tristate
rlabel metal2 s 4324 0 4380 800 6 wbs_dat_o[8]
port 596 nsew default tristate
rlabel metal2 s 4692 0 4748 800 6 wbs_dat_o[9]
port 597 nsew default tristate
rlabel metal2 s 1012 0 1068 800 6 wbs_sel_i[0]
port 598 nsew default input
rlabel metal2 s 1564 0 1620 800 6 wbs_sel_i[1]
port 599 nsew default input
rlabel metal2 s 2024 0 2080 800 6 wbs_sel_i[2]
port 600 nsew default input
rlabel metal2 s 2484 0 2540 800 6 wbs_sel_i[3]
port 601 nsew default input
rlabel metal2 s 460 0 516 800 6 wbs_stb_i
port 602 nsew default input
rlabel metal2 s 552 0 608 800 6 wbs_we_i
port 603 nsew default input
rlabel metal4 s 4190 2128 4510 57712 6 VPWR
port 604 nsew default input
rlabel metal4 s 19550 2128 19870 57712 6 VGND
port 605 nsew default input
<< properties >>
string FIXED_BBOX 0 0 59856 60000
<< end >>
