VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX8
  CLASS CORE ;
  FOREIGN INVX8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.320 2.230 0.610 2.310 ;
        RECT 2.160 2.230 2.450 2.310 ;
        RECT 4.000 2.230 4.290 2.310 ;
        RECT 0.320 2.090 4.290 2.230 ;
        RECT 0.320 2.020 0.610 2.090 ;
        RECT 2.160 2.020 2.450 2.090 ;
        RECT 4.000 2.020 4.290 2.090 ;
        RECT 0.390 0.690 0.530 2.020 ;
        RECT 4.070 0.690 4.210 2.020 ;
        RECT 0.320 0.610 0.610 0.690 ;
        RECT 2.160 0.610 2.450 0.690 ;
        RECT 0.320 0.470 2.450 0.610 ;
        RECT 0.320 0.400 0.610 0.470 ;
        RECT 2.160 0.400 2.450 0.470 ;
        RECT 4.000 0.400 4.290 0.690 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.780 1.690 1.070 1.770 ;
        RECT 1.700 1.690 1.990 1.770 ;
        RECT 2.620 1.690 2.910 1.770 ;
        RECT 3.540 1.690 3.830 1.770 ;
        RECT 0.780 1.550 3.830 1.690 ;
        RECT 0.780 1.480 1.070 1.550 ;
        RECT 1.700 1.480 1.990 1.550 ;
        RECT 2.620 1.480 2.910 1.550 ;
        RECT 3.540 1.480 3.830 1.550 ;
        RECT 0.850 1.230 0.990 1.480 ;
        RECT 1.770 1.230 1.910 1.480 ;
        RECT 2.690 1.230 2.830 1.480 ;
        RECT 3.610 1.230 3.750 1.480 ;
        RECT 0.780 0.940 1.070 1.230 ;
        RECT 1.700 0.940 1.990 1.230 ;
        RECT 2.620 0.940 2.910 1.230 ;
        RECT 3.540 0.940 3.830 1.230 ;
    END
  END A
END INVX8
END LIBRARY

