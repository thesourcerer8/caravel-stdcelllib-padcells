VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1145.470 89.660 1145.790 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 1145.470 89.520 2899.310 89.660 ;
        RECT 1145.470 89.460 1145.790 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 1145.500 89.460 1145.760 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 1150.920 1996.210 1151.200 2000.000 ;
        RECT 1145.560 1996.070 1151.200 1996.210 ;
        RECT 1145.560 89.750 1145.700 1996.070 ;
        RECT 1150.920 1996.000 1151.200 1996.070 ;
        RECT 1145.500 89.430 1145.760 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1234.250 2429.200 1234.570 2429.260 ;
        RECT 2900.830 2429.200 2901.150 2429.260 ;
        RECT 1234.250 2429.060 2901.150 2429.200 ;
        RECT 1234.250 2429.000 1234.570 2429.060 ;
        RECT 2900.830 2429.000 2901.150 2429.060 ;
        RECT 1229.650 2009.300 1229.970 2009.360 ;
        RECT 1234.250 2009.300 1234.570 2009.360 ;
        RECT 1229.650 2009.160 1234.570 2009.300 ;
        RECT 1229.650 2009.100 1229.970 2009.160 ;
        RECT 1234.250 2009.100 1234.570 2009.160 ;
      LAYER via ;
        RECT 1234.280 2429.000 1234.540 2429.260 ;
        RECT 2900.860 2429.000 2901.120 2429.260 ;
        RECT 1229.680 2009.100 1229.940 2009.360 ;
        RECT 1234.280 2009.100 1234.540 2009.360 ;
      LAYER met2 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
        RECT 2900.920 2429.290 2901.060 2433.875 ;
        RECT 1234.280 2428.970 1234.540 2429.290 ;
        RECT 2900.860 2428.970 2901.120 2429.290 ;
        RECT 1234.340 2009.390 1234.480 2428.970 ;
        RECT 1229.680 2009.070 1229.940 2009.390 ;
        RECT 1234.280 2009.070 1234.540 2009.390 ;
        RECT 1229.740 2000.000 1229.880 2009.070 ;
        RECT 1229.580 1999.540 1229.880 2000.000 ;
        RECT 1229.580 1996.000 1229.860 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1241.150 2663.800 1241.470 2663.860 ;
        RECT 2900.830 2663.800 2901.150 2663.860 ;
        RECT 1241.150 2663.660 2901.150 2663.800 ;
        RECT 1241.150 2663.600 1241.470 2663.660 ;
        RECT 2900.830 2663.600 2901.150 2663.660 ;
      LAYER via ;
        RECT 1241.180 2663.600 1241.440 2663.860 ;
        RECT 2900.860 2663.600 2901.120 2663.860 ;
      LAYER met2 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
        RECT 2900.920 2663.890 2901.060 2669.155 ;
        RECT 1241.180 2663.570 1241.440 2663.890 ;
        RECT 2900.860 2663.570 2901.120 2663.890 ;
        RECT 1241.240 2000.290 1241.380 2663.570 ;
        RECT 1239.400 2000.150 1241.380 2000.290 ;
        RECT 1237.400 1999.610 1237.680 2000.000 ;
        RECT 1239.400 1999.610 1239.540 2000.150 ;
        RECT 1237.400 1999.470 1239.540 1999.610 ;
        RECT 1237.400 1996.000 1237.680 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
      LAYER met3 ;
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1248.050 2898.400 1248.370 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 1248.050 2898.260 2901.150 2898.400 ;
        RECT 1248.050 2898.200 1248.370 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
      LAYER via ;
        RECT 1248.080 2898.200 1248.340 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 1248.080 2898.170 1248.340 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 1248.140 2001.650 1248.280 2898.170 ;
        RECT 1247.680 2001.510 1248.280 2001.650 ;
        RECT 1245.220 1999.610 1245.500 2000.000 ;
        RECT 1247.680 1999.610 1247.820 2001.510 ;
        RECT 1245.220 1999.470 1247.820 1999.610 ;
        RECT 1245.220 1996.000 1245.500 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1255.410 3133.000 1255.730 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 1255.410 3132.860 2901.150 3133.000 ;
        RECT 1255.410 3132.800 1255.730 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
      LAYER via ;
        RECT 1255.440 3132.800 1255.700 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 1255.440 3132.770 1255.700 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 1253.500 1999.610 1253.780 2000.000 ;
        RECT 1255.500 1999.610 1255.640 3132.770 ;
        RECT 1253.500 1999.470 1255.640 1999.610 ;
        RECT 1253.500 1996.000 1253.780 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1262.310 3367.600 1262.630 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 1262.310 3367.460 2901.150 3367.600 ;
        RECT 1262.310 3367.400 1262.630 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
      LAYER via ;
        RECT 1262.340 3367.400 1262.600 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 1262.340 3367.370 1262.600 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 1261.320 1999.610 1261.600 2000.000 ;
        RECT 1262.400 1999.610 1262.540 3367.370 ;
        RECT 1261.320 1999.470 1262.540 1999.610 ;
        RECT 1261.320 1996.000 1261.600 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1269.210 3501.560 1269.530 3501.620 ;
        RECT 2798.250 3501.560 2798.570 3501.620 ;
        RECT 1269.210 3501.420 2798.570 3501.560 ;
        RECT 1269.210 3501.360 1269.530 3501.420 ;
        RECT 2798.250 3501.360 2798.570 3501.420 ;
      LAYER via ;
        RECT 1269.240 3501.360 1269.500 3501.620 ;
        RECT 2798.280 3501.360 2798.540 3501.620 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.650 2798.480 3517.600 ;
        RECT 1269.240 3501.330 1269.500 3501.650 ;
        RECT 2798.280 3501.330 2798.540 3501.650 ;
        RECT 1269.300 2000.000 1269.440 3501.330 ;
        RECT 1269.140 1999.540 1269.440 2000.000 ;
        RECT 1269.140 1996.000 1269.420 1999.540 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1283.010 3502.920 1283.330 3502.980 ;
        RECT 2473.950 3502.920 2474.270 3502.980 ;
        RECT 1283.010 3502.780 2474.270 3502.920 ;
        RECT 1283.010 3502.720 1283.330 3502.780 ;
        RECT 2473.950 3502.720 2474.270 3502.780 ;
        RECT 1277.030 2010.660 1277.350 2010.720 ;
        RECT 1283.010 2010.660 1283.330 2010.720 ;
        RECT 1277.030 2010.520 1283.330 2010.660 ;
        RECT 1277.030 2010.460 1277.350 2010.520 ;
        RECT 1283.010 2010.460 1283.330 2010.520 ;
      LAYER via ;
        RECT 1283.040 3502.720 1283.300 3502.980 ;
        RECT 2473.980 3502.720 2474.240 3502.980 ;
        RECT 1277.060 2010.460 1277.320 2010.720 ;
        RECT 1283.040 2010.460 1283.300 2010.720 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3503.010 2474.180 3517.600 ;
        RECT 1283.040 3502.690 1283.300 3503.010 ;
        RECT 2473.980 3502.690 2474.240 3503.010 ;
        RECT 1283.100 2010.750 1283.240 3502.690 ;
        RECT 1277.060 2010.430 1277.320 2010.750 ;
        RECT 1283.040 2010.430 1283.300 2010.750 ;
        RECT 1277.120 2000.000 1277.260 2010.430 ;
        RECT 1276.960 1999.540 1277.260 2000.000 ;
        RECT 1276.960 1996.000 1277.240 1999.540 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1289.910 3504.280 1290.230 3504.340 ;
        RECT 2149.190 3504.280 2149.510 3504.340 ;
        RECT 1289.910 3504.140 2149.510 3504.280 ;
        RECT 1289.910 3504.080 1290.230 3504.140 ;
        RECT 2149.190 3504.080 2149.510 3504.140 ;
        RECT 1284.850 2010.660 1285.170 2010.720 ;
        RECT 1289.910 2010.660 1290.230 2010.720 ;
        RECT 1284.850 2010.520 1290.230 2010.660 ;
        RECT 1284.850 2010.460 1285.170 2010.520 ;
        RECT 1289.910 2010.460 1290.230 2010.520 ;
      LAYER via ;
        RECT 1289.940 3504.080 1290.200 3504.340 ;
        RECT 2149.220 3504.080 2149.480 3504.340 ;
        RECT 1284.880 2010.460 1285.140 2010.720 ;
        RECT 1289.940 2010.460 1290.200 2010.720 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3504.370 2149.420 3517.600 ;
        RECT 1289.940 3504.050 1290.200 3504.370 ;
        RECT 2149.220 3504.050 2149.480 3504.370 ;
        RECT 1290.000 2010.750 1290.140 3504.050 ;
        RECT 1284.880 2010.430 1285.140 2010.750 ;
        RECT 1289.940 2010.430 1290.200 2010.750 ;
        RECT 1284.940 2000.000 1285.080 2010.430 ;
        RECT 1284.780 1999.540 1285.080 2000.000 ;
        RECT 1284.780 1996.000 1285.060 1999.540 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1296.810 3500.880 1297.130 3500.940 ;
        RECT 1824.890 3500.880 1825.210 3500.940 ;
        RECT 1296.810 3500.740 1825.210 3500.880 ;
        RECT 1296.810 3500.680 1297.130 3500.740 ;
        RECT 1824.890 3500.680 1825.210 3500.740 ;
        RECT 1292.670 2010.320 1292.990 2010.380 ;
        RECT 1296.810 2010.320 1297.130 2010.380 ;
        RECT 1292.670 2010.180 1297.130 2010.320 ;
        RECT 1292.670 2010.120 1292.990 2010.180 ;
        RECT 1296.810 2010.120 1297.130 2010.180 ;
      LAYER via ;
        RECT 1296.840 3500.680 1297.100 3500.940 ;
        RECT 1824.920 3500.680 1825.180 3500.940 ;
        RECT 1292.700 2010.120 1292.960 2010.380 ;
        RECT 1296.840 2010.120 1297.100 2010.380 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3500.970 1825.120 3517.600 ;
        RECT 1296.840 3500.650 1297.100 3500.970 ;
        RECT 1824.920 3500.650 1825.180 3500.970 ;
        RECT 1296.900 2010.410 1297.040 3500.650 ;
        RECT 1292.700 2010.090 1292.960 2010.410 ;
        RECT 1296.840 2010.090 1297.100 2010.410 ;
        RECT 1292.760 2000.000 1292.900 2010.090 ;
        RECT 1292.600 1999.540 1292.900 2000.000 ;
        RECT 1292.600 1996.000 1292.880 1999.540 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1499.285 3332.765 1499.455 3422.355 ;
        RECT 1498.365 3008.405 1498.535 3042.915 ;
        RECT 1499.285 2946.525 1499.455 2994.635 ;
        RECT 1498.365 2428.705 1498.535 2463.215 ;
        RECT 1498.365 2331.805 1498.535 2366.655 ;
        RECT 1497.445 2201.245 1497.615 2249.355 ;
        RECT 1497.905 2138.685 1498.075 2184.075 ;
        RECT 1498.365 2028.525 1498.535 2076.975 ;
        RECT 1309.305 2010.505 1309.475 2013.055 ;
      LAYER mcon ;
        RECT 1499.285 3422.185 1499.455 3422.355 ;
        RECT 1498.365 3042.745 1498.535 3042.915 ;
        RECT 1499.285 2994.465 1499.455 2994.635 ;
        RECT 1498.365 2463.045 1498.535 2463.215 ;
        RECT 1498.365 2366.485 1498.535 2366.655 ;
        RECT 1497.445 2249.185 1497.615 2249.355 ;
        RECT 1497.905 2183.905 1498.075 2184.075 ;
        RECT 1498.365 2076.805 1498.535 2076.975 ;
        RECT 1309.305 2012.885 1309.475 2013.055 ;
      LAYER met1 ;
        RECT 1498.290 3443.080 1498.610 3443.140 ;
        RECT 1500.590 3443.080 1500.910 3443.140 ;
        RECT 1498.290 3442.940 1500.910 3443.080 ;
        RECT 1498.290 3442.880 1498.610 3442.940 ;
        RECT 1500.590 3442.880 1500.910 3442.940 ;
        RECT 1497.830 3422.340 1498.150 3422.400 ;
        RECT 1499.225 3422.340 1499.515 3422.385 ;
        RECT 1497.830 3422.200 1499.515 3422.340 ;
        RECT 1497.830 3422.140 1498.150 3422.200 ;
        RECT 1499.225 3422.155 1499.515 3422.200 ;
        RECT 1499.225 3332.920 1499.515 3332.965 ;
        RECT 1499.670 3332.920 1499.990 3332.980 ;
        RECT 1499.225 3332.780 1499.990 3332.920 ;
        RECT 1499.225 3332.735 1499.515 3332.780 ;
        RECT 1499.670 3332.720 1499.990 3332.780 ;
        RECT 1498.290 3236.360 1498.610 3236.420 ;
        RECT 1498.750 3236.360 1499.070 3236.420 ;
        RECT 1498.290 3236.220 1499.070 3236.360 ;
        RECT 1498.290 3236.160 1498.610 3236.220 ;
        RECT 1498.750 3236.160 1499.070 3236.220 ;
        RECT 1498.290 3202.020 1498.610 3202.080 ;
        RECT 1498.750 3202.020 1499.070 3202.080 ;
        RECT 1498.290 3201.880 1499.070 3202.020 ;
        RECT 1498.290 3201.820 1498.610 3201.880 ;
        RECT 1498.750 3201.820 1499.070 3201.880 ;
        RECT 1497.830 3153.400 1498.150 3153.460 ;
        RECT 1498.750 3153.400 1499.070 3153.460 ;
        RECT 1497.830 3153.260 1499.070 3153.400 ;
        RECT 1497.830 3153.200 1498.150 3153.260 ;
        RECT 1498.750 3153.200 1499.070 3153.260 ;
        RECT 1497.830 3056.840 1498.150 3056.900 ;
        RECT 1498.750 3056.840 1499.070 3056.900 ;
        RECT 1497.830 3056.700 1499.070 3056.840 ;
        RECT 1497.830 3056.640 1498.150 3056.700 ;
        RECT 1498.750 3056.640 1499.070 3056.700 ;
        RECT 1498.290 3042.900 1498.610 3042.960 ;
        RECT 1498.095 3042.760 1498.610 3042.900 ;
        RECT 1498.290 3042.700 1498.610 3042.760 ;
        RECT 1498.305 3008.560 1498.595 3008.605 ;
        RECT 1499.210 3008.560 1499.530 3008.620 ;
        RECT 1498.305 3008.420 1499.530 3008.560 ;
        RECT 1498.305 3008.375 1498.595 3008.420 ;
        RECT 1499.210 3008.360 1499.530 3008.420 ;
        RECT 1499.210 2994.620 1499.530 2994.680 ;
        RECT 1499.015 2994.480 1499.530 2994.620 ;
        RECT 1499.210 2994.420 1499.530 2994.480 ;
        RECT 1499.225 2946.680 1499.515 2946.725 ;
        RECT 1499.670 2946.680 1499.990 2946.740 ;
        RECT 1499.225 2946.540 1499.990 2946.680 ;
        RECT 1499.225 2946.495 1499.515 2946.540 ;
        RECT 1499.670 2946.480 1499.990 2946.540 ;
        RECT 1499.670 2912.340 1499.990 2912.400 ;
        RECT 1499.300 2912.200 1499.990 2912.340 ;
        RECT 1499.300 2911.720 1499.440 2912.200 ;
        RECT 1499.670 2912.140 1499.990 2912.200 ;
        RECT 1499.210 2911.460 1499.530 2911.720 ;
        RECT 1497.830 2815.580 1498.150 2815.840 ;
        RECT 1497.920 2815.160 1498.060 2815.580 ;
        RECT 1497.830 2814.900 1498.150 2815.160 ;
        RECT 1497.830 2767.500 1498.150 2767.560 ;
        RECT 1497.460 2767.360 1498.150 2767.500 ;
        RECT 1497.460 2766.880 1497.600 2767.360 ;
        RECT 1497.830 2767.300 1498.150 2767.360 ;
        RECT 1497.370 2766.620 1497.690 2766.880 ;
        RECT 1496.450 2718.540 1496.770 2718.600 ;
        RECT 1497.370 2718.540 1497.690 2718.600 ;
        RECT 1496.450 2718.400 1497.690 2718.540 ;
        RECT 1496.450 2718.340 1496.770 2718.400 ;
        RECT 1497.370 2718.340 1497.690 2718.400 ;
        RECT 1497.830 2656.660 1498.150 2656.720 ;
        RECT 1498.750 2656.660 1499.070 2656.720 ;
        RECT 1497.830 2656.520 1499.070 2656.660 ;
        RECT 1497.830 2656.460 1498.150 2656.520 ;
        RECT 1498.750 2656.460 1499.070 2656.520 ;
        RECT 1498.750 2622.120 1499.070 2622.380 ;
        RECT 1498.840 2621.980 1498.980 2622.120 ;
        RECT 1499.210 2621.980 1499.530 2622.040 ;
        RECT 1498.840 2621.840 1499.530 2621.980 ;
        RECT 1499.210 2621.780 1499.530 2621.840 ;
        RECT 1498.290 2560.100 1498.610 2560.160 ;
        RECT 1499.670 2560.100 1499.990 2560.160 ;
        RECT 1498.290 2559.960 1499.990 2560.100 ;
        RECT 1498.290 2559.900 1498.610 2559.960 ;
        RECT 1499.670 2559.900 1499.990 2559.960 ;
        RECT 1498.750 2511.820 1499.070 2511.880 ;
        RECT 1499.670 2511.820 1499.990 2511.880 ;
        RECT 1498.750 2511.680 1499.990 2511.820 ;
        RECT 1498.750 2511.620 1499.070 2511.680 ;
        RECT 1499.670 2511.620 1499.990 2511.680 ;
        RECT 1498.290 2463.200 1498.610 2463.260 ;
        RECT 1498.095 2463.060 1498.610 2463.200 ;
        RECT 1498.290 2463.000 1498.610 2463.060 ;
        RECT 1498.290 2428.860 1498.610 2428.920 ;
        RECT 1498.095 2428.720 1498.610 2428.860 ;
        RECT 1498.290 2428.660 1498.610 2428.720 ;
        RECT 1497.830 2380.580 1498.150 2380.640 ;
        RECT 1498.750 2380.580 1499.070 2380.640 ;
        RECT 1497.830 2380.440 1499.070 2380.580 ;
        RECT 1497.830 2380.380 1498.150 2380.440 ;
        RECT 1498.750 2380.380 1499.070 2380.440 ;
        RECT 1498.290 2366.640 1498.610 2366.700 ;
        RECT 1498.095 2366.500 1498.610 2366.640 ;
        RECT 1498.290 2366.440 1498.610 2366.500 ;
        RECT 1498.290 2331.960 1498.610 2332.020 ;
        RECT 1498.095 2331.820 1498.610 2331.960 ;
        RECT 1498.290 2331.760 1498.610 2331.820 ;
        RECT 1496.910 2304.420 1497.230 2304.480 ;
        RECT 1498.750 2304.420 1499.070 2304.480 ;
        RECT 1496.910 2304.280 1499.070 2304.420 ;
        RECT 1496.910 2304.220 1497.230 2304.280 ;
        RECT 1498.750 2304.220 1499.070 2304.280 ;
        RECT 1497.370 2249.340 1497.690 2249.400 ;
        RECT 1497.175 2249.200 1497.690 2249.340 ;
        RECT 1497.370 2249.140 1497.690 2249.200 ;
        RECT 1497.385 2201.400 1497.675 2201.445 ;
        RECT 1497.830 2201.400 1498.150 2201.460 ;
        RECT 1497.385 2201.260 1498.150 2201.400 ;
        RECT 1497.385 2201.215 1497.675 2201.260 ;
        RECT 1497.830 2201.200 1498.150 2201.260 ;
        RECT 1497.830 2184.060 1498.150 2184.120 ;
        RECT 1497.635 2183.920 1498.150 2184.060 ;
        RECT 1497.830 2183.860 1498.150 2183.920 ;
        RECT 1497.830 2138.840 1498.150 2138.900 ;
        RECT 1497.635 2138.700 1498.150 2138.840 ;
        RECT 1497.830 2138.640 1498.150 2138.700 ;
        RECT 1498.305 2076.960 1498.595 2077.005 ;
        RECT 1498.750 2076.960 1499.070 2077.020 ;
        RECT 1498.305 2076.820 1499.070 2076.960 ;
        RECT 1498.305 2076.775 1498.595 2076.820 ;
        RECT 1498.750 2076.760 1499.070 2076.820 ;
        RECT 1498.290 2028.680 1498.610 2028.740 ;
        RECT 1498.095 2028.540 1498.610 2028.680 ;
        RECT 1498.290 2028.480 1498.610 2028.540 ;
        RECT 1300.950 2013.040 1301.270 2013.100 ;
        RECT 1309.245 2013.040 1309.535 2013.085 ;
        RECT 1300.950 2012.900 1309.535 2013.040 ;
        RECT 1300.950 2012.840 1301.270 2012.900 ;
        RECT 1309.245 2012.855 1309.535 2012.900 ;
        RECT 1309.245 2010.660 1309.535 2010.705 ;
        RECT 1498.290 2010.660 1498.610 2010.720 ;
        RECT 1309.245 2010.520 1498.610 2010.660 ;
        RECT 1309.245 2010.475 1309.535 2010.520 ;
        RECT 1498.290 2010.460 1498.610 2010.520 ;
      LAYER via ;
        RECT 1498.320 3442.880 1498.580 3443.140 ;
        RECT 1500.620 3442.880 1500.880 3443.140 ;
        RECT 1497.860 3422.140 1498.120 3422.400 ;
        RECT 1499.700 3332.720 1499.960 3332.980 ;
        RECT 1498.320 3236.160 1498.580 3236.420 ;
        RECT 1498.780 3236.160 1499.040 3236.420 ;
        RECT 1498.320 3201.820 1498.580 3202.080 ;
        RECT 1498.780 3201.820 1499.040 3202.080 ;
        RECT 1497.860 3153.200 1498.120 3153.460 ;
        RECT 1498.780 3153.200 1499.040 3153.460 ;
        RECT 1497.860 3056.640 1498.120 3056.900 ;
        RECT 1498.780 3056.640 1499.040 3056.900 ;
        RECT 1498.320 3042.700 1498.580 3042.960 ;
        RECT 1499.240 3008.360 1499.500 3008.620 ;
        RECT 1499.240 2994.420 1499.500 2994.680 ;
        RECT 1499.700 2946.480 1499.960 2946.740 ;
        RECT 1499.700 2912.140 1499.960 2912.400 ;
        RECT 1499.240 2911.460 1499.500 2911.720 ;
        RECT 1497.860 2815.580 1498.120 2815.840 ;
        RECT 1497.860 2814.900 1498.120 2815.160 ;
        RECT 1497.860 2767.300 1498.120 2767.560 ;
        RECT 1497.400 2766.620 1497.660 2766.880 ;
        RECT 1496.480 2718.340 1496.740 2718.600 ;
        RECT 1497.400 2718.340 1497.660 2718.600 ;
        RECT 1497.860 2656.460 1498.120 2656.720 ;
        RECT 1498.780 2656.460 1499.040 2656.720 ;
        RECT 1498.780 2622.120 1499.040 2622.380 ;
        RECT 1499.240 2621.780 1499.500 2622.040 ;
        RECT 1498.320 2559.900 1498.580 2560.160 ;
        RECT 1499.700 2559.900 1499.960 2560.160 ;
        RECT 1498.780 2511.620 1499.040 2511.880 ;
        RECT 1499.700 2511.620 1499.960 2511.880 ;
        RECT 1498.320 2463.000 1498.580 2463.260 ;
        RECT 1498.320 2428.660 1498.580 2428.920 ;
        RECT 1497.860 2380.380 1498.120 2380.640 ;
        RECT 1498.780 2380.380 1499.040 2380.640 ;
        RECT 1498.320 2366.440 1498.580 2366.700 ;
        RECT 1498.320 2331.760 1498.580 2332.020 ;
        RECT 1496.940 2304.220 1497.200 2304.480 ;
        RECT 1498.780 2304.220 1499.040 2304.480 ;
        RECT 1497.400 2249.140 1497.660 2249.400 ;
        RECT 1497.860 2201.200 1498.120 2201.460 ;
        RECT 1497.860 2183.860 1498.120 2184.120 ;
        RECT 1497.860 2138.640 1498.120 2138.900 ;
        RECT 1498.780 2076.760 1499.040 2077.020 ;
        RECT 1498.320 2028.480 1498.580 2028.740 ;
        RECT 1300.980 2012.840 1301.240 2013.100 ;
        RECT 1498.320 2010.460 1498.580 2010.720 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3443.170 1500.820 3517.600 ;
        RECT 1498.320 3442.850 1498.580 3443.170 ;
        RECT 1500.620 3442.850 1500.880 3443.170 ;
        RECT 1498.380 3429.650 1498.520 3442.850 ;
        RECT 1497.920 3429.510 1498.520 3429.650 ;
        RECT 1497.920 3422.430 1498.060 3429.510 ;
        RECT 1497.860 3422.110 1498.120 3422.430 ;
        RECT 1499.700 3332.690 1499.960 3333.010 ;
        RECT 1499.760 3298.410 1499.900 3332.690 ;
        RECT 1498.840 3298.270 1499.900 3298.410 ;
        RECT 1498.840 3236.450 1498.980 3298.270 ;
        RECT 1498.320 3236.130 1498.580 3236.450 ;
        RECT 1498.780 3236.130 1499.040 3236.450 ;
        RECT 1498.380 3202.110 1498.520 3236.130 ;
        RECT 1498.320 3201.790 1498.580 3202.110 ;
        RECT 1498.780 3201.790 1499.040 3202.110 ;
        RECT 1498.840 3153.490 1498.980 3201.790 ;
        RECT 1497.860 3153.170 1498.120 3153.490 ;
        RECT 1498.780 3153.170 1499.040 3153.490 ;
        RECT 1497.920 3152.890 1498.060 3153.170 ;
        RECT 1497.920 3152.750 1498.520 3152.890 ;
        RECT 1498.380 3105.290 1498.520 3152.750 ;
        RECT 1498.380 3105.150 1498.980 3105.290 ;
        RECT 1498.840 3056.930 1498.980 3105.150 ;
        RECT 1497.860 3056.610 1498.120 3056.930 ;
        RECT 1498.780 3056.610 1499.040 3056.930 ;
        RECT 1497.920 3056.330 1498.060 3056.610 ;
        RECT 1497.920 3056.190 1498.520 3056.330 ;
        RECT 1498.380 3042.990 1498.520 3056.190 ;
        RECT 1498.320 3042.670 1498.580 3042.990 ;
        RECT 1499.240 3008.330 1499.500 3008.650 ;
        RECT 1499.300 2994.710 1499.440 3008.330 ;
        RECT 1499.240 2994.390 1499.500 2994.710 ;
        RECT 1499.700 2946.450 1499.960 2946.770 ;
        RECT 1499.760 2912.430 1499.900 2946.450 ;
        RECT 1499.700 2912.110 1499.960 2912.430 ;
        RECT 1499.240 2911.430 1499.500 2911.750 ;
        RECT 1499.300 2863.210 1499.440 2911.430 ;
        RECT 1498.380 2863.070 1499.440 2863.210 ;
        RECT 1498.380 2849.610 1498.520 2863.070 ;
        RECT 1497.920 2849.470 1498.520 2849.610 ;
        RECT 1497.920 2815.870 1498.060 2849.470 ;
        RECT 1497.860 2815.550 1498.120 2815.870 ;
        RECT 1497.860 2814.870 1498.120 2815.190 ;
        RECT 1497.920 2802.805 1498.060 2814.870 ;
        RECT 1497.850 2802.435 1498.130 2802.805 ;
        RECT 1497.850 2801.755 1498.130 2802.125 ;
        RECT 1497.920 2767.590 1498.060 2801.755 ;
        RECT 1497.860 2767.270 1498.120 2767.590 ;
        RECT 1497.400 2766.590 1497.660 2766.910 ;
        RECT 1497.460 2746.365 1497.600 2766.590 ;
        RECT 1496.470 2745.995 1496.750 2746.365 ;
        RECT 1497.390 2745.995 1497.670 2746.365 ;
        RECT 1496.540 2718.630 1496.680 2745.995 ;
        RECT 1496.480 2718.310 1496.740 2718.630 ;
        RECT 1497.400 2718.310 1497.660 2718.630 ;
        RECT 1497.460 2697.970 1497.600 2718.310 ;
        RECT 1497.460 2697.830 1498.060 2697.970 ;
        RECT 1497.920 2656.750 1498.060 2697.830 ;
        RECT 1497.860 2656.430 1498.120 2656.750 ;
        RECT 1498.780 2656.430 1499.040 2656.750 ;
        RECT 1498.840 2622.410 1498.980 2656.430 ;
        RECT 1498.780 2622.090 1499.040 2622.410 ;
        RECT 1499.240 2621.750 1499.500 2622.070 ;
        RECT 1499.300 2608.325 1499.440 2621.750 ;
        RECT 1498.310 2607.955 1498.590 2608.325 ;
        RECT 1499.230 2607.955 1499.510 2608.325 ;
        RECT 1498.380 2560.190 1498.520 2607.955 ;
        RECT 1498.320 2559.870 1498.580 2560.190 ;
        RECT 1499.700 2559.870 1499.960 2560.190 ;
        RECT 1499.760 2511.910 1499.900 2559.870 ;
        RECT 1498.780 2511.765 1499.040 2511.910 ;
        RECT 1497.390 2511.395 1497.670 2511.765 ;
        RECT 1498.770 2511.395 1499.050 2511.765 ;
        RECT 1499.700 2511.590 1499.960 2511.910 ;
        RECT 1497.460 2463.485 1497.600 2511.395 ;
        RECT 1497.390 2463.115 1497.670 2463.485 ;
        RECT 1498.310 2463.115 1498.590 2463.485 ;
        RECT 1498.320 2462.970 1498.580 2463.115 ;
        RECT 1498.320 2428.630 1498.580 2428.950 ;
        RECT 1498.380 2415.090 1498.520 2428.630 ;
        RECT 1498.380 2414.950 1498.980 2415.090 ;
        RECT 1498.840 2380.670 1498.980 2414.950 ;
        RECT 1497.860 2380.410 1498.120 2380.670 ;
        RECT 1497.860 2380.350 1498.520 2380.410 ;
        RECT 1498.780 2380.350 1499.040 2380.670 ;
        RECT 1497.920 2380.270 1498.520 2380.350 ;
        RECT 1498.380 2366.730 1498.520 2380.270 ;
        RECT 1498.320 2366.410 1498.580 2366.730 ;
        RECT 1498.320 2331.730 1498.580 2332.050 ;
        RECT 1498.380 2318.530 1498.520 2331.730 ;
        RECT 1498.380 2318.390 1498.980 2318.530 ;
        RECT 1498.840 2304.510 1498.980 2318.390 ;
        RECT 1496.940 2304.190 1497.200 2304.510 ;
        RECT 1498.780 2304.190 1499.040 2304.510 ;
        RECT 1497.000 2256.650 1497.140 2304.190 ;
        RECT 1497.000 2256.510 1497.600 2256.650 ;
        RECT 1497.460 2249.430 1497.600 2256.510 ;
        RECT 1497.400 2249.110 1497.660 2249.430 ;
        RECT 1497.860 2201.170 1498.120 2201.490 ;
        RECT 1497.920 2184.150 1498.060 2201.170 ;
        RECT 1497.860 2183.830 1498.120 2184.150 ;
        RECT 1497.860 2138.610 1498.120 2138.930 ;
        RECT 1497.920 2090.730 1498.060 2138.610 ;
        RECT 1497.920 2090.590 1498.980 2090.730 ;
        RECT 1498.840 2077.050 1498.980 2090.590 ;
        RECT 1498.780 2076.730 1499.040 2077.050 ;
        RECT 1498.320 2028.450 1498.580 2028.770 ;
        RECT 1300.980 2012.810 1301.240 2013.130 ;
        RECT 1301.040 2000.000 1301.180 2012.810 ;
        RECT 1498.380 2010.750 1498.520 2028.450 ;
        RECT 1498.320 2010.430 1498.580 2010.750 ;
        RECT 1300.880 1999.540 1301.180 2000.000 ;
        RECT 1300.880 1996.000 1301.160 1999.540 ;
      LAYER via2 ;
        RECT 1497.850 2802.480 1498.130 2802.760 ;
        RECT 1497.850 2801.800 1498.130 2802.080 ;
        RECT 1496.470 2746.040 1496.750 2746.320 ;
        RECT 1497.390 2746.040 1497.670 2746.320 ;
        RECT 1498.310 2608.000 1498.590 2608.280 ;
        RECT 1499.230 2608.000 1499.510 2608.280 ;
        RECT 1497.390 2511.440 1497.670 2511.720 ;
        RECT 1498.770 2511.440 1499.050 2511.720 ;
        RECT 1497.390 2463.160 1497.670 2463.440 ;
        RECT 1498.310 2463.160 1498.590 2463.440 ;
      LAYER met3 ;
        RECT 1497.825 2802.770 1498.155 2802.785 ;
        RECT 1497.150 2802.470 1498.155 2802.770 ;
        RECT 1497.150 2802.090 1497.450 2802.470 ;
        RECT 1497.825 2802.455 1498.155 2802.470 ;
        RECT 1497.825 2802.090 1498.155 2802.105 ;
        RECT 1497.150 2801.790 1498.155 2802.090 ;
        RECT 1497.825 2801.775 1498.155 2801.790 ;
        RECT 1496.445 2746.330 1496.775 2746.345 ;
        RECT 1497.365 2746.330 1497.695 2746.345 ;
        RECT 1496.445 2746.030 1497.695 2746.330 ;
        RECT 1496.445 2746.015 1496.775 2746.030 ;
        RECT 1497.365 2746.015 1497.695 2746.030 ;
        RECT 1498.285 2608.290 1498.615 2608.305 ;
        RECT 1499.205 2608.290 1499.535 2608.305 ;
        RECT 1498.285 2607.990 1499.535 2608.290 ;
        RECT 1498.285 2607.975 1498.615 2607.990 ;
        RECT 1499.205 2607.975 1499.535 2607.990 ;
        RECT 1497.365 2511.730 1497.695 2511.745 ;
        RECT 1498.745 2511.730 1499.075 2511.745 ;
        RECT 1497.365 2511.430 1499.075 2511.730 ;
        RECT 1497.365 2511.415 1497.695 2511.430 ;
        RECT 1498.745 2511.415 1499.075 2511.430 ;
        RECT 1497.365 2463.450 1497.695 2463.465 ;
        RECT 1498.285 2463.450 1498.615 2463.465 ;
        RECT 1497.365 2463.150 1498.615 2463.450 ;
        RECT 1497.365 2463.135 1497.695 2463.150 ;
        RECT 1498.285 2463.135 1498.615 2463.150 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1158.810 2004.540 1159.130 2004.600 ;
        RECT 1472.990 2004.540 1473.310 2004.600 ;
        RECT 1158.810 2004.400 1473.310 2004.540 ;
        RECT 1158.810 2004.340 1159.130 2004.400 ;
        RECT 1472.990 2004.340 1473.310 2004.400 ;
        RECT 1472.990 324.260 1473.310 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 1472.990 324.120 2899.310 324.260 ;
        RECT 1472.990 324.060 1473.310 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 1158.840 2004.340 1159.100 2004.600 ;
        RECT 1473.020 2004.340 1473.280 2004.600 ;
        RECT 1473.020 324.060 1473.280 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 1158.840 2004.310 1159.100 2004.630 ;
        RECT 1473.020 2004.310 1473.280 2004.630 ;
        RECT 1158.900 2000.000 1159.040 2004.310 ;
        RECT 1158.740 1999.540 1159.040 2000.000 ;
        RECT 1158.740 1996.000 1159.020 1999.540 ;
        RECT 1473.080 324.350 1473.220 2004.310 ;
        RECT 1473.020 324.030 1473.280 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
        RECT 1308.770 2010.660 1309.090 2010.720 ;
        RECT 1292.300 2010.520 1309.090 2010.660 ;
        RECT 1179.510 2010.320 1179.830 2010.380 ;
        RECT 1292.300 2010.320 1292.440 2010.520 ;
        RECT 1308.770 2010.460 1309.090 2010.520 ;
        RECT 1179.510 2010.180 1292.440 2010.320 ;
        RECT 1179.510 2010.120 1179.830 2010.180 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
        RECT 1179.540 2010.120 1179.800 2010.380 ;
        RECT 1308.800 2010.460 1309.060 2010.720 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 2010.410 1179.740 3498.270 ;
        RECT 1308.800 2010.430 1309.060 2010.750 ;
        RECT 1179.540 2010.090 1179.800 2010.410 ;
        RECT 1308.860 2000.000 1309.000 2010.430 ;
        RECT 1308.700 1999.540 1309.000 2000.000 ;
        RECT 1308.700 1996.000 1308.980 1999.540 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3498.500 851.850 3498.560 ;
        RECT 855.210 3498.500 855.530 3498.560 ;
        RECT 851.530 3498.360 855.530 3498.500 ;
        RECT 851.530 3498.300 851.850 3498.360 ;
        RECT 855.210 3498.300 855.530 3498.360 ;
        RECT 855.210 2014.740 855.530 2014.800 ;
        RECT 1316.590 2014.740 1316.910 2014.800 ;
        RECT 855.210 2014.600 1316.910 2014.740 ;
        RECT 855.210 2014.540 855.530 2014.600 ;
        RECT 1316.590 2014.540 1316.910 2014.600 ;
      LAYER via ;
        RECT 851.560 3498.300 851.820 3498.560 ;
        RECT 855.240 3498.300 855.500 3498.560 ;
        RECT 855.240 2014.540 855.500 2014.800 ;
        RECT 1316.620 2014.540 1316.880 2014.800 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3498.590 851.760 3517.600 ;
        RECT 851.560 3498.270 851.820 3498.590 ;
        RECT 855.240 3498.270 855.500 3498.590 ;
        RECT 855.300 2014.830 855.440 3498.270 ;
        RECT 855.240 2014.510 855.500 2014.830 ;
        RECT 1316.620 2014.510 1316.880 2014.830 ;
        RECT 1316.680 2000.000 1316.820 2014.510 ;
        RECT 1316.520 1999.540 1316.820 2000.000 ;
        RECT 1316.520 1996.000 1316.800 1999.540 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 530.910 3498.500 531.230 3498.560 ;
        RECT 527.230 3498.360 531.230 3498.500 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 530.910 3498.300 531.230 3498.360 ;
        RECT 530.910 2014.060 531.230 2014.120 ;
        RECT 530.910 2013.920 1291.980 2014.060 ;
        RECT 530.910 2013.860 531.230 2013.920 ;
        RECT 1291.840 2013.720 1291.980 2013.920 ;
        RECT 1324.410 2013.720 1324.730 2013.780 ;
        RECT 1291.840 2013.580 1324.730 2013.720 ;
        RECT 1324.410 2013.520 1324.730 2013.580 ;
      LAYER via ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 530.940 3498.300 531.200 3498.560 ;
        RECT 530.940 2013.860 531.200 2014.120 ;
        RECT 1324.440 2013.520 1324.700 2013.780 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 530.940 3498.270 531.200 3498.590 ;
        RECT 531.000 2014.150 531.140 3498.270 ;
        RECT 530.940 2013.830 531.200 2014.150 ;
        RECT 1324.440 2013.490 1324.700 2013.810 ;
        RECT 1324.500 2000.000 1324.640 2013.490 ;
        RECT 1324.340 1999.540 1324.640 2000.000 ;
        RECT 1324.340 1996.000 1324.620 1999.540 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1300.565 2012.885 1300.735 2014.075 ;
        RECT 1311.145 2012.885 1311.315 2014.075 ;
      LAYER mcon ;
        RECT 1300.565 2013.905 1300.735 2014.075 ;
        RECT 1311.145 2013.905 1311.315 2014.075 ;
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 206.610 3501.900 206.930 3501.960 ;
        RECT 202.470 3501.760 206.930 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 206.610 3501.700 206.930 3501.760 ;
        RECT 1300.505 2014.060 1300.795 2014.105 ;
        RECT 1311.085 2014.060 1311.375 2014.105 ;
        RECT 1300.505 2013.920 1311.375 2014.060 ;
        RECT 1300.505 2013.875 1300.795 2013.920 ;
        RECT 1311.085 2013.875 1311.375 2013.920 ;
        RECT 206.610 2013.380 206.930 2013.440 ;
        RECT 206.610 2013.240 1291.060 2013.380 ;
        RECT 206.610 2013.180 206.930 2013.240 ;
        RECT 1290.920 2013.040 1291.060 2013.240 ;
        RECT 1300.505 2013.040 1300.795 2013.085 ;
        RECT 1290.920 2012.900 1300.795 2013.040 ;
        RECT 1300.505 2012.855 1300.795 2012.900 ;
        RECT 1311.085 2013.040 1311.375 2013.085 ;
        RECT 1332.230 2013.040 1332.550 2013.100 ;
        RECT 1311.085 2012.900 1332.550 2013.040 ;
        RECT 1311.085 2012.855 1311.375 2012.900 ;
        RECT 1332.230 2012.840 1332.550 2012.900 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 206.640 3501.700 206.900 3501.960 ;
        RECT 206.640 2013.180 206.900 2013.440 ;
        RECT 1332.260 2012.840 1332.520 2013.100 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 206.640 3501.670 206.900 3501.990 ;
        RECT 206.700 2013.470 206.840 3501.670 ;
        RECT 206.640 2013.150 206.900 2013.470 ;
        RECT 1332.260 2012.810 1332.520 2013.130 ;
        RECT 1332.320 2000.000 1332.460 2012.810 ;
        RECT 1332.160 1999.540 1332.460 2000.000 ;
        RECT 1332.160 1996.000 1332.440 1999.540 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1313.905 2010.165 1314.075 2012.715 ;
      LAYER mcon ;
        RECT 1313.905 2012.545 1314.075 2012.715 ;
      LAYER met1 ;
        RECT 17.090 2012.700 17.410 2012.760 ;
        RECT 1313.845 2012.700 1314.135 2012.745 ;
        RECT 17.090 2012.560 1314.135 2012.700 ;
        RECT 17.090 2012.500 17.410 2012.560 ;
        RECT 1313.845 2012.515 1314.135 2012.560 ;
        RECT 1313.845 2010.320 1314.135 2010.365 ;
        RECT 1340.050 2010.320 1340.370 2010.380 ;
        RECT 1313.845 2010.180 1340.370 2010.320 ;
        RECT 1313.845 2010.135 1314.135 2010.180 ;
        RECT 1340.050 2010.120 1340.370 2010.180 ;
      LAYER via ;
        RECT 17.120 2012.500 17.380 2012.760 ;
        RECT 1340.080 2010.120 1340.340 2010.380 ;
      LAYER met2 ;
        RECT 17.110 3411.035 17.390 3411.405 ;
        RECT 17.180 2012.790 17.320 3411.035 ;
        RECT 17.120 2012.470 17.380 2012.790 ;
        RECT 1340.080 2010.090 1340.340 2010.410 ;
        RECT 1340.140 2000.000 1340.280 2010.090 ;
        RECT 1339.980 1999.540 1340.280 2000.000 ;
        RECT 1339.980 1996.000 1340.260 1999.540 ;
      LAYER via2 ;
        RECT 17.110 3411.080 17.390 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.085 3411.370 17.415 3411.385 ;
        RECT -4.800 3411.070 17.415 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.085 3411.055 17.415 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1305.625 2012.205 1305.795 2015.095 ;
      LAYER mcon ;
        RECT 1305.625 2014.925 1305.795 2015.095 ;
      LAYER met1 ;
        RECT 1305.565 2015.080 1305.855 2015.125 ;
        RECT 1305.565 2014.940 1317.280 2015.080 ;
        RECT 1305.565 2014.895 1305.855 2014.940 ;
        RECT 1317.140 2014.740 1317.280 2014.940 ;
        RECT 1346.030 2014.740 1346.350 2014.800 ;
        RECT 1317.140 2014.600 1346.350 2014.740 ;
        RECT 1346.030 2014.540 1346.350 2014.600 ;
        RECT 17.550 2012.360 17.870 2012.420 ;
        RECT 1305.565 2012.360 1305.855 2012.405 ;
        RECT 17.550 2012.220 1305.855 2012.360 ;
        RECT 17.550 2012.160 17.870 2012.220 ;
        RECT 1305.565 2012.175 1305.855 2012.220 ;
      LAYER via ;
        RECT 1346.060 2014.540 1346.320 2014.800 ;
        RECT 17.580 2012.160 17.840 2012.420 ;
      LAYER met2 ;
        RECT 17.570 3124.075 17.850 3124.445 ;
        RECT 17.640 2012.450 17.780 3124.075 ;
        RECT 1346.060 2014.510 1346.320 2014.830 ;
        RECT 17.580 2012.130 17.840 2012.450 ;
        RECT 1346.120 1999.610 1346.260 2014.510 ;
        RECT 1347.800 1999.610 1348.080 2000.000 ;
        RECT 1346.120 1999.470 1348.080 1999.610 ;
        RECT 1347.800 1996.000 1348.080 1999.470 ;
      LAYER via2 ;
        RECT 17.570 3124.120 17.850 3124.400 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.545 3124.410 17.875 3124.425 ;
        RECT -4.800 3124.110 17.875 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.545 3124.095 17.875 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.470 2012.020 18.790 2012.080 ;
        RECT 1356.150 2012.020 1356.470 2012.080 ;
        RECT 18.470 2011.880 1356.470 2012.020 ;
        RECT 18.470 2011.820 18.790 2011.880 ;
        RECT 1356.150 2011.820 1356.470 2011.880 ;
      LAYER via ;
        RECT 18.500 2011.820 18.760 2012.080 ;
        RECT 1356.180 2011.820 1356.440 2012.080 ;
      LAYER met2 ;
        RECT 18.490 2836.435 18.770 2836.805 ;
        RECT 18.560 2012.110 18.700 2836.435 ;
        RECT 18.500 2011.790 18.760 2012.110 ;
        RECT 1356.180 2011.790 1356.440 2012.110 ;
        RECT 1356.240 2000.000 1356.380 2011.790 ;
        RECT 1356.080 1999.540 1356.380 2000.000 ;
        RECT 1356.080 1996.000 1356.360 1999.540 ;
      LAYER via2 ;
        RECT 18.490 2836.480 18.770 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 18.465 2836.770 18.795 2836.785 ;
        RECT -4.800 2836.470 18.795 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 18.465 2836.455 18.795 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.390 2011.680 19.710 2011.740 ;
        RECT 1363.970 2011.680 1364.290 2011.740 ;
        RECT 19.390 2011.540 1364.290 2011.680 ;
        RECT 19.390 2011.480 19.710 2011.540 ;
        RECT 1363.970 2011.480 1364.290 2011.540 ;
      LAYER via ;
        RECT 19.420 2011.480 19.680 2011.740 ;
        RECT 1364.000 2011.480 1364.260 2011.740 ;
      LAYER met2 ;
        RECT 19.410 2549.475 19.690 2549.845 ;
        RECT 19.480 2011.770 19.620 2549.475 ;
        RECT 19.420 2011.450 19.680 2011.770 ;
        RECT 1364.000 2011.450 1364.260 2011.770 ;
        RECT 1364.060 2000.000 1364.200 2011.450 ;
        RECT 1363.900 1999.540 1364.200 2000.000 ;
        RECT 1363.900 1996.000 1364.180 1999.540 ;
      LAYER via2 ;
        RECT 19.410 2549.520 19.690 2549.800 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 19.385 2549.810 19.715 2549.825 ;
        RECT -4.800 2549.510 19.715 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 19.385 2549.495 19.715 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 2011.340 20.630 2011.400 ;
        RECT 1371.790 2011.340 1372.110 2011.400 ;
        RECT 20.310 2011.200 1372.110 2011.340 ;
        RECT 20.310 2011.140 20.630 2011.200 ;
        RECT 1371.790 2011.140 1372.110 2011.200 ;
      LAYER via ;
        RECT 20.340 2011.140 20.600 2011.400 ;
        RECT 1371.820 2011.140 1372.080 2011.400 ;
      LAYER met2 ;
        RECT 20.330 2261.835 20.610 2262.205 ;
        RECT 20.400 2011.430 20.540 2261.835 ;
        RECT 20.340 2011.110 20.600 2011.430 ;
        RECT 1371.820 2011.110 1372.080 2011.430 ;
        RECT 1371.880 2000.000 1372.020 2011.110 ;
        RECT 1371.720 1999.540 1372.020 2000.000 ;
        RECT 1371.720 1996.000 1372.000 1999.540 ;
      LAYER via2 ;
        RECT 20.330 2261.880 20.610 2262.160 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 20.305 2262.170 20.635 2262.185 ;
        RECT -4.800 2261.870 20.635 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 20.305 2261.855 20.635 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 54.810 1999.780 55.130 1999.840 ;
        RECT 1378.230 1999.780 1378.550 1999.840 ;
        RECT 54.810 1999.640 1378.550 1999.780 ;
        RECT 54.810 1999.580 55.130 1999.640 ;
        RECT 1378.230 1999.580 1378.550 1999.640 ;
        RECT 15.710 1980.060 16.030 1980.120 ;
        RECT 54.810 1980.060 55.130 1980.120 ;
        RECT 15.710 1979.920 55.130 1980.060 ;
        RECT 15.710 1979.860 16.030 1979.920 ;
        RECT 54.810 1979.860 55.130 1979.920 ;
      LAYER via ;
        RECT 54.840 1999.580 55.100 1999.840 ;
        RECT 1378.260 1999.580 1378.520 1999.840 ;
        RECT 15.740 1979.860 16.000 1980.120 ;
        RECT 54.840 1979.860 55.100 1980.120 ;
      LAYER met2 ;
        RECT 54.840 1999.550 55.100 1999.870 ;
        RECT 1378.260 1999.610 1378.520 1999.870 ;
        RECT 1379.540 1999.610 1379.820 2000.000 ;
        RECT 1378.260 1999.550 1379.820 1999.610 ;
        RECT 54.900 1980.150 55.040 1999.550 ;
        RECT 1378.320 1999.470 1379.820 1999.550 ;
        RECT 1379.540 1996.000 1379.820 1999.470 ;
        RECT 15.740 1979.830 16.000 1980.150 ;
        RECT 54.840 1979.830 55.100 1980.150 ;
        RECT 15.800 1975.245 15.940 1979.830 ;
        RECT 15.730 1974.875 16.010 1975.245 ;
      LAYER via2 ;
        RECT 15.730 1974.920 16.010 1975.200 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 15.705 1975.210 16.035 1975.225 ;
        RECT -4.800 1974.910 16.035 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 15.705 1974.895 16.035 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1168.010 1998.420 1168.330 1998.480 ;
        RECT 1459.650 1998.420 1459.970 1998.480 ;
        RECT 1168.010 1998.280 1459.970 1998.420 ;
        RECT 1168.010 1998.220 1168.330 1998.280 ;
        RECT 1459.650 1998.220 1459.970 1998.280 ;
        RECT 1459.650 558.860 1459.970 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 1459.650 558.720 2899.310 558.860 ;
        RECT 1459.650 558.660 1459.970 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 1168.040 1998.220 1168.300 1998.480 ;
        RECT 1459.680 1998.220 1459.940 1998.480 ;
        RECT 1459.680 558.660 1459.940 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 1166.560 1998.250 1166.840 2000.000 ;
        RECT 1168.040 1998.250 1168.300 1998.510 ;
        RECT 1166.560 1998.190 1168.300 1998.250 ;
        RECT 1459.680 1998.190 1459.940 1998.510 ;
        RECT 1166.560 1998.110 1168.240 1998.190 ;
        RECT 1166.560 1996.000 1166.840 1998.110 ;
        RECT 1459.740 558.950 1459.880 1998.190 ;
        RECT 1459.680 558.630 1459.940 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 65.390 2006.580 65.710 2006.640 ;
        RECT 1387.430 2006.580 1387.750 2006.640 ;
        RECT 65.390 2006.440 1387.750 2006.580 ;
        RECT 65.390 2006.380 65.710 2006.440 ;
        RECT 1387.430 2006.380 1387.750 2006.440 ;
        RECT 17.090 1690.380 17.410 1690.440 ;
        RECT 65.390 1690.380 65.710 1690.440 ;
        RECT 17.090 1690.240 65.710 1690.380 ;
        RECT 17.090 1690.180 17.410 1690.240 ;
        RECT 65.390 1690.180 65.710 1690.240 ;
      LAYER via ;
        RECT 65.420 2006.380 65.680 2006.640 ;
        RECT 1387.460 2006.380 1387.720 2006.640 ;
        RECT 17.120 1690.180 17.380 1690.440 ;
        RECT 65.420 1690.180 65.680 1690.440 ;
      LAYER met2 ;
        RECT 65.420 2006.350 65.680 2006.670 ;
        RECT 1387.460 2006.350 1387.720 2006.670 ;
        RECT 65.480 1690.470 65.620 2006.350 ;
        RECT 1387.520 2000.000 1387.660 2006.350 ;
        RECT 1387.360 1999.540 1387.660 2000.000 ;
        RECT 1387.360 1996.000 1387.640 1999.540 ;
        RECT 17.120 1690.150 17.380 1690.470 ;
        RECT 65.420 1690.150 65.680 1690.470 ;
        RECT 17.180 1687.605 17.320 1690.150 ;
        RECT 17.110 1687.235 17.390 1687.605 ;
      LAYER via2 ;
        RECT 17.110 1687.280 17.390 1687.560 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 17.085 1687.570 17.415 1687.585 ;
        RECT -4.800 1687.270 17.415 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 17.085 1687.255 17.415 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1135.810 1999.100 1136.130 1999.160 ;
        RECT 1393.870 1999.100 1394.190 1999.160 ;
        RECT 1135.810 1998.960 1394.190 1999.100 ;
        RECT 1135.810 1998.900 1136.130 1998.960 ;
        RECT 1393.870 1998.900 1394.190 1998.960 ;
        RECT 15.250 1476.520 15.570 1476.580 ;
        RECT 1135.810 1476.520 1136.130 1476.580 ;
        RECT 15.250 1476.380 1136.130 1476.520 ;
        RECT 15.250 1476.320 15.570 1476.380 ;
        RECT 1135.810 1476.320 1136.130 1476.380 ;
      LAYER via ;
        RECT 1135.840 1998.900 1136.100 1999.160 ;
        RECT 1393.900 1998.900 1394.160 1999.160 ;
        RECT 15.280 1476.320 15.540 1476.580 ;
        RECT 1135.840 1476.320 1136.100 1476.580 ;
      LAYER met2 ;
        RECT 1135.840 1998.870 1136.100 1999.190 ;
        RECT 1393.900 1998.930 1394.160 1999.190 ;
        RECT 1395.180 1998.930 1395.460 2000.000 ;
        RECT 1393.900 1998.870 1395.460 1998.930 ;
        RECT 1135.900 1476.610 1136.040 1998.870 ;
        RECT 1393.960 1998.790 1395.460 1998.870 ;
        RECT 1395.180 1996.000 1395.460 1998.790 ;
        RECT 15.280 1476.290 15.540 1476.610 ;
        RECT 1135.840 1476.290 1136.100 1476.610 ;
        RECT 15.340 1472.045 15.480 1476.290 ;
        RECT 15.270 1471.675 15.550 1472.045 ;
      LAYER via2 ;
        RECT 15.270 1471.720 15.550 1472.000 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 15.245 1472.010 15.575 1472.025 ;
        RECT -4.800 1471.710 15.575 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 15.245 1471.695 15.575 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1128.910 2005.560 1129.230 2005.620 ;
        RECT 1403.530 2005.560 1403.850 2005.620 ;
        RECT 1128.910 2005.420 1403.850 2005.560 ;
        RECT 1128.910 2005.360 1129.230 2005.420 ;
        RECT 1403.530 2005.360 1403.850 2005.420 ;
        RECT 17.090 1262.660 17.410 1262.720 ;
        RECT 1128.910 1262.660 1129.230 1262.720 ;
        RECT 17.090 1262.520 1129.230 1262.660 ;
        RECT 17.090 1262.460 17.410 1262.520 ;
        RECT 1128.910 1262.460 1129.230 1262.520 ;
      LAYER via ;
        RECT 1128.940 2005.360 1129.200 2005.620 ;
        RECT 1403.560 2005.360 1403.820 2005.620 ;
        RECT 17.120 1262.460 17.380 1262.720 ;
        RECT 1128.940 1262.460 1129.200 1262.720 ;
      LAYER met2 ;
        RECT 1128.940 2005.330 1129.200 2005.650 ;
        RECT 1403.560 2005.330 1403.820 2005.650 ;
        RECT 1129.000 1262.750 1129.140 2005.330 ;
        RECT 1403.620 2000.000 1403.760 2005.330 ;
        RECT 1403.460 1999.540 1403.760 2000.000 ;
        RECT 1403.460 1996.000 1403.740 1999.540 ;
        RECT 17.120 1262.430 17.380 1262.750 ;
        RECT 1128.940 1262.430 1129.200 1262.750 ;
        RECT 17.180 1256.485 17.320 1262.430 ;
        RECT 17.110 1256.115 17.390 1256.485 ;
      LAYER via2 ;
        RECT 17.110 1256.160 17.390 1256.440 ;
      LAYER met3 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 17.085 1256.450 17.415 1256.465 ;
        RECT -4.800 1256.150 17.415 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 17.085 1256.135 17.415 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1114.650 1998.760 1114.970 1998.820 ;
        RECT 1409.510 1998.760 1409.830 1998.820 ;
        RECT 1114.650 1998.620 1409.830 1998.760 ;
        RECT 1114.650 1998.560 1114.970 1998.620 ;
        RECT 1409.510 1998.560 1409.830 1998.620 ;
        RECT 17.090 1041.660 17.410 1041.720 ;
        RECT 1114.650 1041.660 1114.970 1041.720 ;
        RECT 17.090 1041.520 1114.970 1041.660 ;
        RECT 17.090 1041.460 17.410 1041.520 ;
        RECT 1114.650 1041.460 1114.970 1041.520 ;
      LAYER via ;
        RECT 1114.680 1998.560 1114.940 1998.820 ;
        RECT 1409.540 1998.560 1409.800 1998.820 ;
        RECT 17.120 1041.460 17.380 1041.720 ;
        RECT 1114.680 1041.460 1114.940 1041.720 ;
      LAYER met2 ;
        RECT 1411.280 1998.930 1411.560 2000.000 ;
        RECT 1409.600 1998.850 1411.560 1998.930 ;
        RECT 1114.680 1998.530 1114.940 1998.850 ;
        RECT 1409.540 1998.790 1411.560 1998.850 ;
        RECT 1409.540 1998.530 1409.800 1998.790 ;
        RECT 1114.740 1041.750 1114.880 1998.530 ;
        RECT 1411.280 1996.000 1411.560 1998.790 ;
        RECT 17.120 1041.430 17.380 1041.750 ;
        RECT 1114.680 1041.430 1114.940 1041.750 ;
        RECT 17.180 1040.925 17.320 1041.430 ;
        RECT 17.110 1040.555 17.390 1040.925 ;
      LAYER via2 ;
        RECT 17.110 1040.600 17.390 1040.880 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 17.085 1040.890 17.415 1040.905 ;
        RECT -4.800 1040.590 17.415 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 17.085 1040.575 17.415 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1093.490 2003.860 1093.810 2003.920 ;
        RECT 1419.170 2003.860 1419.490 2003.920 ;
        RECT 1093.490 2003.720 1419.490 2003.860 ;
        RECT 1093.490 2003.660 1093.810 2003.720 ;
        RECT 1419.170 2003.660 1419.490 2003.720 ;
        RECT 17.550 827.800 17.870 827.860 ;
        RECT 1093.490 827.800 1093.810 827.860 ;
        RECT 17.550 827.660 1093.810 827.800 ;
        RECT 17.550 827.600 17.870 827.660 ;
        RECT 1093.490 827.600 1093.810 827.660 ;
      LAYER via ;
        RECT 1093.520 2003.660 1093.780 2003.920 ;
        RECT 1419.200 2003.660 1419.460 2003.920 ;
        RECT 17.580 827.600 17.840 827.860 ;
        RECT 1093.520 827.600 1093.780 827.860 ;
      LAYER met2 ;
        RECT 1093.520 2003.630 1093.780 2003.950 ;
        RECT 1419.200 2003.630 1419.460 2003.950 ;
        RECT 1093.580 827.890 1093.720 2003.630 ;
        RECT 1419.260 2000.000 1419.400 2003.630 ;
        RECT 1419.100 1999.540 1419.400 2000.000 ;
        RECT 1419.100 1996.000 1419.380 1999.540 ;
        RECT 17.580 827.570 17.840 827.890 ;
        RECT 1093.520 827.570 1093.780 827.890 ;
        RECT 17.640 825.365 17.780 827.570 ;
        RECT 17.570 824.995 17.850 825.365 ;
      LAYER via2 ;
        RECT 17.570 825.040 17.850 825.320 ;
      LAYER met3 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 17.545 825.330 17.875 825.345 ;
        RECT -4.800 825.030 17.875 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 17.545 825.015 17.875 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1079.690 1997.060 1080.010 1997.120 ;
        RECT 1425.150 1997.060 1425.470 1997.120 ;
        RECT 1079.690 1996.920 1425.470 1997.060 ;
        RECT 1079.690 1996.860 1080.010 1996.920 ;
        RECT 1425.150 1996.860 1425.470 1996.920 ;
        RECT 17.090 613.940 17.410 614.000 ;
        RECT 1079.690 613.940 1080.010 614.000 ;
        RECT 17.090 613.800 1080.010 613.940 ;
        RECT 17.090 613.740 17.410 613.800 ;
        RECT 1079.690 613.740 1080.010 613.800 ;
      LAYER via ;
        RECT 1079.720 1996.860 1079.980 1997.120 ;
        RECT 1425.180 1996.860 1425.440 1997.120 ;
        RECT 17.120 613.740 17.380 614.000 ;
        RECT 1079.720 613.740 1079.980 614.000 ;
      LAYER met2 ;
        RECT 1079.720 1996.830 1079.980 1997.150 ;
        RECT 1425.180 1996.890 1425.440 1997.150 ;
        RECT 1426.920 1996.890 1427.200 2000.000 ;
        RECT 1425.180 1996.830 1427.200 1996.890 ;
        RECT 1079.780 614.030 1079.920 1996.830 ;
        RECT 1425.240 1996.750 1427.200 1996.830 ;
        RECT 1426.920 1996.000 1427.200 1996.750 ;
        RECT 17.120 613.710 17.380 614.030 ;
        RECT 1079.720 613.710 1079.980 614.030 ;
        RECT 17.180 610.485 17.320 613.710 ;
        RECT 17.110 610.115 17.390 610.485 ;
      LAYER via2 ;
        RECT 17.110 610.160 17.390 610.440 ;
      LAYER met3 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 17.085 610.450 17.415 610.465 ;
        RECT -4.800 610.150 17.415 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 17.085 610.135 17.415 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1072.790 2003.180 1073.110 2003.240 ;
        RECT 1434.810 2003.180 1435.130 2003.240 ;
        RECT 1072.790 2003.040 1435.130 2003.180 ;
        RECT 1072.790 2002.980 1073.110 2003.040 ;
        RECT 1434.810 2002.980 1435.130 2003.040 ;
        RECT 17.090 400.080 17.410 400.140 ;
        RECT 1072.790 400.080 1073.110 400.140 ;
        RECT 17.090 399.940 1073.110 400.080 ;
        RECT 17.090 399.880 17.410 399.940 ;
        RECT 1072.790 399.880 1073.110 399.940 ;
      LAYER via ;
        RECT 1072.820 2002.980 1073.080 2003.240 ;
        RECT 1434.840 2002.980 1435.100 2003.240 ;
        RECT 17.120 399.880 17.380 400.140 ;
        RECT 1072.820 399.880 1073.080 400.140 ;
      LAYER met2 ;
        RECT 1072.820 2002.950 1073.080 2003.270 ;
        RECT 1434.840 2002.950 1435.100 2003.270 ;
        RECT 1072.880 400.170 1073.020 2002.950 ;
        RECT 1434.900 2000.000 1435.040 2002.950 ;
        RECT 1434.740 1999.540 1435.040 2000.000 ;
        RECT 1434.740 1996.000 1435.020 1999.540 ;
        RECT 17.120 399.850 17.380 400.170 ;
        RECT 1072.820 399.850 1073.080 400.170 ;
        RECT 17.180 394.925 17.320 399.850 ;
        RECT 17.110 394.555 17.390 394.925 ;
      LAYER via2 ;
        RECT 17.110 394.600 17.390 394.880 ;
      LAYER met3 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 17.085 394.890 17.415 394.905 ;
        RECT -4.800 394.590 17.415 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 17.085 394.575 17.415 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1441.785 1995.885 1441.955 1996.735 ;
      LAYER mcon ;
        RECT 1441.785 1996.565 1441.955 1996.735 ;
      LAYER met1 ;
        RECT 1441.710 1996.720 1442.030 1996.780 ;
        RECT 1441.515 1996.580 1442.030 1996.720 ;
        RECT 1441.710 1996.520 1442.030 1996.580 ;
        RECT 1065.890 1996.040 1066.210 1996.100 ;
        RECT 1441.725 1996.040 1442.015 1996.085 ;
        RECT 1065.890 1995.900 1442.015 1996.040 ;
        RECT 1065.890 1995.840 1066.210 1995.900 ;
        RECT 1441.725 1995.855 1442.015 1995.900 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 1065.890 179.420 1066.210 179.480 ;
        RECT 17.090 179.280 1066.210 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 1065.890 179.220 1066.210 179.280 ;
      LAYER via ;
        RECT 1441.740 1996.520 1442.000 1996.780 ;
        RECT 1065.920 1995.840 1066.180 1996.100 ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 1065.920 179.220 1066.180 179.480 ;
      LAYER met2 ;
        RECT 1442.560 1996.890 1442.840 2000.000 ;
        RECT 1441.800 1996.810 1442.840 1996.890 ;
        RECT 1441.740 1996.750 1442.840 1996.810 ;
        RECT 1441.740 1996.490 1442.000 1996.750 ;
        RECT 1065.920 1995.810 1066.180 1996.130 ;
        RECT 1442.560 1996.000 1442.840 1996.750 ;
        RECT 1065.980 179.510 1066.120 1995.810 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 1065.920 179.190 1066.180 179.510 ;
      LAYER via2 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.085 179.015 17.415 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1174.450 2004.880 1174.770 2004.940 ;
        RECT 1487.250 2004.880 1487.570 2004.940 ;
        RECT 1174.450 2004.740 1487.570 2004.880 ;
        RECT 1174.450 2004.680 1174.770 2004.740 ;
        RECT 1487.250 2004.680 1487.570 2004.740 ;
        RECT 1487.250 793.460 1487.570 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 1487.250 793.320 2899.310 793.460 ;
        RECT 1487.250 793.260 1487.570 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 1174.480 2004.680 1174.740 2004.940 ;
        RECT 1487.280 2004.680 1487.540 2004.940 ;
        RECT 1487.280 793.260 1487.540 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 1174.480 2004.650 1174.740 2004.970 ;
        RECT 1487.280 2004.650 1487.540 2004.970 ;
        RECT 1174.540 2000.000 1174.680 2004.650 ;
        RECT 1174.380 1999.540 1174.680 2000.000 ;
        RECT 1174.380 1996.000 1174.660 1999.540 ;
        RECT 1487.340 793.550 1487.480 2004.650 ;
        RECT 1487.280 793.230 1487.540 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
        RECT 2898.985 792.010 2899.315 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1183.650 1998.080 1183.970 1998.140 ;
        RECT 1494.150 1998.080 1494.470 1998.140 ;
        RECT 1183.650 1997.940 1494.470 1998.080 ;
        RECT 1183.650 1997.880 1183.970 1997.940 ;
        RECT 1494.150 1997.880 1494.470 1997.940 ;
        RECT 1494.150 1028.060 1494.470 1028.120 ;
        RECT 2898.990 1028.060 2899.310 1028.120 ;
        RECT 1494.150 1027.920 2899.310 1028.060 ;
        RECT 1494.150 1027.860 1494.470 1027.920 ;
        RECT 2898.990 1027.860 2899.310 1027.920 ;
      LAYER via ;
        RECT 1183.680 1997.880 1183.940 1998.140 ;
        RECT 1494.180 1997.880 1494.440 1998.140 ;
        RECT 1494.180 1027.860 1494.440 1028.120 ;
        RECT 2899.020 1027.860 2899.280 1028.120 ;
      LAYER met2 ;
        RECT 1182.200 1998.250 1182.480 2000.000 ;
        RECT 1182.200 1998.170 1183.880 1998.250 ;
        RECT 1182.200 1998.110 1183.940 1998.170 ;
        RECT 1182.200 1996.000 1182.480 1998.110 ;
        RECT 1183.680 1997.850 1183.940 1998.110 ;
        RECT 1494.180 1997.850 1494.440 1998.170 ;
        RECT 1494.240 1028.150 1494.380 1997.850 ;
        RECT 1494.180 1027.830 1494.440 1028.150 ;
        RECT 2899.020 1027.830 2899.280 1028.150 ;
        RECT 2899.080 1026.645 2899.220 1027.830 ;
        RECT 2899.010 1026.275 2899.290 1026.645 ;
      LAYER via2 ;
        RECT 2899.010 1026.320 2899.290 1026.600 ;
      LAYER met3 ;
        RECT 2898.985 1026.610 2899.315 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2898.985 1026.310 2924.800 1026.610 ;
        RECT 2898.985 1026.295 2899.315 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1190.090 2004.200 1190.410 2004.260 ;
        RECT 1507.950 2004.200 1508.270 2004.260 ;
        RECT 1190.090 2004.060 1508.270 2004.200 ;
        RECT 1190.090 2004.000 1190.410 2004.060 ;
        RECT 1507.950 2004.000 1508.270 2004.060 ;
        RECT 1507.950 1262.660 1508.270 1262.720 ;
        RECT 2898.990 1262.660 2899.310 1262.720 ;
        RECT 1507.950 1262.520 2899.310 1262.660 ;
        RECT 1507.950 1262.460 1508.270 1262.520 ;
        RECT 2898.990 1262.460 2899.310 1262.520 ;
      LAYER via ;
        RECT 1190.120 2004.000 1190.380 2004.260 ;
        RECT 1507.980 2004.000 1508.240 2004.260 ;
        RECT 1507.980 1262.460 1508.240 1262.720 ;
        RECT 2899.020 1262.460 2899.280 1262.720 ;
      LAYER met2 ;
        RECT 1190.120 2003.970 1190.380 2004.290 ;
        RECT 1507.980 2003.970 1508.240 2004.290 ;
        RECT 1190.180 2000.000 1190.320 2003.970 ;
        RECT 1190.020 1999.540 1190.320 2000.000 ;
        RECT 1190.020 1996.000 1190.300 1999.540 ;
        RECT 1508.040 1262.750 1508.180 2003.970 ;
        RECT 1507.980 1262.430 1508.240 1262.750 ;
        RECT 2899.020 1262.430 2899.280 1262.750 ;
        RECT 2899.080 1261.245 2899.220 1262.430 ;
        RECT 2899.010 1260.875 2899.290 1261.245 ;
      LAYER via2 ;
        RECT 2899.010 1260.920 2899.290 1261.200 ;
      LAYER met3 ;
        RECT 2898.985 1261.210 2899.315 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2898.985 1260.910 2924.800 1261.210 ;
        RECT 2898.985 1260.895 2899.315 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1199.290 1997.400 1199.610 1997.460 ;
        RECT 1514.850 1997.400 1515.170 1997.460 ;
        RECT 1199.290 1997.260 1515.170 1997.400 ;
        RECT 1199.290 1997.200 1199.610 1997.260 ;
        RECT 1514.850 1997.200 1515.170 1997.260 ;
        RECT 1514.850 1497.260 1515.170 1497.320 ;
        RECT 2898.990 1497.260 2899.310 1497.320 ;
        RECT 1514.850 1497.120 2899.310 1497.260 ;
        RECT 1514.850 1497.060 1515.170 1497.120 ;
        RECT 2898.990 1497.060 2899.310 1497.120 ;
      LAYER via ;
        RECT 1199.320 1997.200 1199.580 1997.460 ;
        RECT 1514.880 1997.200 1515.140 1997.460 ;
        RECT 1514.880 1497.060 1515.140 1497.320 ;
        RECT 2899.020 1497.060 2899.280 1497.320 ;
      LAYER met2 ;
        RECT 1197.840 1997.570 1198.120 2000.000 ;
        RECT 1197.840 1997.490 1199.520 1997.570 ;
        RECT 1197.840 1997.430 1199.580 1997.490 ;
        RECT 1197.840 1996.000 1198.120 1997.430 ;
        RECT 1199.320 1997.170 1199.580 1997.430 ;
        RECT 1514.880 1997.170 1515.140 1997.490 ;
        RECT 1514.940 1497.350 1515.080 1997.170 ;
        RECT 1514.880 1497.030 1515.140 1497.350 ;
        RECT 2899.020 1497.030 2899.280 1497.350 ;
        RECT 2899.080 1495.845 2899.220 1497.030 ;
        RECT 2899.010 1495.475 2899.290 1495.845 ;
      LAYER via2 ;
        RECT 2899.010 1495.520 2899.290 1495.800 ;
      LAYER met3 ;
        RECT 2898.985 1495.810 2899.315 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2898.985 1495.510 2924.800 1495.810 ;
        RECT 2898.985 1495.495 2899.315 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1206.190 2005.900 1206.510 2005.960 ;
        RECT 1452.290 2005.900 1452.610 2005.960 ;
        RECT 1206.190 2005.760 1452.610 2005.900 ;
        RECT 1206.190 2005.700 1206.510 2005.760 ;
        RECT 1452.290 2005.700 1452.610 2005.760 ;
        RECT 1452.290 1731.860 1452.610 1731.920 ;
        RECT 2898.990 1731.860 2899.310 1731.920 ;
        RECT 1452.290 1731.720 2899.310 1731.860 ;
        RECT 1452.290 1731.660 1452.610 1731.720 ;
        RECT 2898.990 1731.660 2899.310 1731.720 ;
      LAYER via ;
        RECT 1206.220 2005.700 1206.480 2005.960 ;
        RECT 1452.320 2005.700 1452.580 2005.960 ;
        RECT 1452.320 1731.660 1452.580 1731.920 ;
        RECT 2899.020 1731.660 2899.280 1731.920 ;
      LAYER met2 ;
        RECT 1206.220 2005.670 1206.480 2005.990 ;
        RECT 1452.320 2005.670 1452.580 2005.990 ;
        RECT 1206.280 2000.000 1206.420 2005.670 ;
        RECT 1206.120 1999.540 1206.420 2000.000 ;
        RECT 1206.120 1996.000 1206.400 1999.540 ;
        RECT 1452.380 1731.950 1452.520 2005.670 ;
        RECT 1452.320 1731.630 1452.580 1731.950 ;
        RECT 2899.020 1731.630 2899.280 1731.950 ;
        RECT 2899.080 1730.445 2899.220 1731.630 ;
        RECT 2899.010 1730.075 2899.290 1730.445 ;
      LAYER via2 ;
        RECT 2899.010 1730.120 2899.290 1730.400 ;
      LAYER met3 ;
        RECT 2898.985 1730.410 2899.315 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2898.985 1730.110 2924.800 1730.410 ;
        RECT 2898.985 1730.095 2899.315 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1214.470 1999.440 1214.790 1999.500 ;
        RECT 1453.210 1999.440 1453.530 1999.500 ;
        RECT 1214.470 1999.300 1453.530 1999.440 ;
        RECT 1214.470 1999.240 1214.790 1999.300 ;
        RECT 1453.210 1999.240 1453.530 1999.300 ;
        RECT 1453.210 1966.460 1453.530 1966.520 ;
        RECT 2898.990 1966.460 2899.310 1966.520 ;
        RECT 1453.210 1966.320 2899.310 1966.460 ;
        RECT 1453.210 1966.260 1453.530 1966.320 ;
        RECT 2898.990 1966.260 2899.310 1966.320 ;
      LAYER via ;
        RECT 1214.500 1999.240 1214.760 1999.500 ;
        RECT 1453.240 1999.240 1453.500 1999.500 ;
        RECT 1453.240 1966.260 1453.500 1966.520 ;
        RECT 2899.020 1966.260 2899.280 1966.520 ;
      LAYER met2 ;
        RECT 1213.940 1999.610 1214.220 2000.000 ;
        RECT 1213.940 1999.530 1214.700 1999.610 ;
        RECT 1213.940 1999.470 1214.760 1999.530 ;
        RECT 1213.940 1996.000 1214.220 1999.470 ;
        RECT 1214.500 1999.210 1214.760 1999.470 ;
        RECT 1453.240 1999.210 1453.500 1999.530 ;
        RECT 1453.300 1966.550 1453.440 1999.210 ;
        RECT 1453.240 1966.230 1453.500 1966.550 ;
        RECT 2899.020 1966.230 2899.280 1966.550 ;
        RECT 2899.080 1965.045 2899.220 1966.230 ;
        RECT 2899.010 1964.675 2899.290 1965.045 ;
      LAYER via2 ;
        RECT 2899.010 1964.720 2899.290 1965.000 ;
      LAYER met3 ;
        RECT 2898.985 1965.010 2899.315 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2898.985 1964.710 2924.800 1965.010 ;
        RECT 2898.985 1964.695 2899.315 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1226.890 2194.600 1227.210 2194.660 ;
        RECT 2900.830 2194.600 2901.150 2194.660 ;
        RECT 1226.890 2194.460 2901.150 2194.600 ;
        RECT 1226.890 2194.400 1227.210 2194.460 ;
        RECT 2900.830 2194.400 2901.150 2194.460 ;
        RECT 1221.830 2009.300 1222.150 2009.360 ;
        RECT 1226.890 2009.300 1227.210 2009.360 ;
        RECT 1221.830 2009.160 1227.210 2009.300 ;
        RECT 1221.830 2009.100 1222.150 2009.160 ;
        RECT 1226.890 2009.100 1227.210 2009.160 ;
      LAYER via ;
        RECT 1226.920 2194.400 1227.180 2194.660 ;
        RECT 2900.860 2194.400 2901.120 2194.660 ;
        RECT 1221.860 2009.100 1222.120 2009.360 ;
        RECT 1226.920 2009.100 1227.180 2009.360 ;
      LAYER met2 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
        RECT 2900.920 2194.690 2901.060 2199.275 ;
        RECT 1226.920 2194.370 1227.180 2194.690 ;
        RECT 2900.860 2194.370 2901.120 2194.690 ;
        RECT 1226.980 2009.390 1227.120 2194.370 ;
        RECT 1221.860 2009.070 1222.120 2009.390 ;
        RECT 1226.920 2009.070 1227.180 2009.390 ;
        RECT 1221.920 2000.000 1222.060 2009.070 ;
        RECT 1221.760 1999.540 1222.060 2000.000 ;
        RECT 1221.760 1996.000 1222.040 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
      LAYER met3 ;
        RECT 2900.825 2199.610 2901.155 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1153.290 2002.500 1153.610 2002.560 ;
        RECT 1521.290 2002.500 1521.610 2002.560 ;
        RECT 1153.290 2002.360 1521.610 2002.500 ;
        RECT 1153.290 2002.300 1153.610 2002.360 ;
        RECT 1521.290 2002.300 1521.610 2002.360 ;
        RECT 1521.290 206.960 1521.610 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 1521.290 206.820 2901.150 206.960 ;
        RECT 1521.290 206.760 1521.610 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 1153.320 2002.300 1153.580 2002.560 ;
        RECT 1521.320 2002.300 1521.580 2002.560 ;
        RECT 1521.320 206.760 1521.580 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 1153.320 2002.270 1153.580 2002.590 ;
        RECT 1521.320 2002.270 1521.580 2002.590 ;
        RECT 1153.380 2000.000 1153.520 2002.270 ;
        RECT 1153.220 1999.540 1153.520 2000.000 ;
        RECT 1153.220 1996.000 1153.500 1999.540 ;
        RECT 1521.380 207.050 1521.520 2002.270 ;
        RECT 1521.320 206.730 1521.580 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1234.710 2546.500 1235.030 2546.560 ;
        RECT 2900.830 2546.500 2901.150 2546.560 ;
        RECT 1234.710 2546.360 2901.150 2546.500 ;
        RECT 1234.710 2546.300 1235.030 2546.360 ;
        RECT 2900.830 2546.300 2901.150 2546.360 ;
      LAYER via ;
        RECT 1234.740 2546.300 1235.000 2546.560 ;
        RECT 2900.860 2546.300 2901.120 2546.560 ;
      LAYER met2 ;
        RECT 2900.850 2551.515 2901.130 2551.885 ;
        RECT 2900.920 2546.590 2901.060 2551.515 ;
        RECT 1234.740 2546.270 1235.000 2546.590 ;
        RECT 2900.860 2546.270 2901.120 2546.590 ;
        RECT 1232.340 1999.610 1232.620 2000.000 ;
        RECT 1234.800 1999.610 1234.940 2546.270 ;
        RECT 1232.340 1999.470 1234.940 1999.610 ;
        RECT 1232.340 1996.000 1232.620 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 2551.560 2901.130 2551.840 ;
      LAYER met3 ;
        RECT 2900.825 2551.850 2901.155 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2900.825 2551.550 2924.800 2551.850 ;
        RECT 2900.825 2551.535 2901.155 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1241.610 2781.100 1241.930 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 1241.610 2780.960 2901.150 2781.100 ;
        RECT 1241.610 2780.900 1241.930 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
      LAYER via ;
        RECT 1241.640 2780.900 1241.900 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 1241.640 2780.870 1241.900 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 1240.160 1999.610 1240.440 2000.000 ;
        RECT 1241.700 1999.610 1241.840 2780.870 ;
        RECT 1240.160 1999.470 1241.840 1999.610 ;
        RECT 1240.160 1996.000 1240.440 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1248.510 3015.700 1248.830 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 1248.510 3015.560 2901.150 3015.700 ;
        RECT 1248.510 3015.500 1248.830 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
      LAYER via ;
        RECT 1248.540 3015.500 1248.800 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 1248.540 3015.470 1248.800 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 1247.980 1999.610 1248.260 2000.000 ;
        RECT 1248.600 1999.610 1248.740 3015.470 ;
        RECT 1247.980 1999.470 1248.740 1999.610 ;
        RECT 1247.980 1996.000 1248.260 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1261.850 3250.300 1262.170 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 1261.850 3250.160 2901.150 3250.300 ;
        RECT 1261.850 3250.100 1262.170 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
        RECT 1255.870 2010.660 1256.190 2010.720 ;
        RECT 1261.850 2010.660 1262.170 2010.720 ;
        RECT 1255.870 2010.520 1262.170 2010.660 ;
        RECT 1255.870 2010.460 1256.190 2010.520 ;
        RECT 1261.850 2010.460 1262.170 2010.520 ;
      LAYER via ;
        RECT 1261.880 3250.100 1262.140 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
        RECT 1255.900 2010.460 1256.160 2010.720 ;
        RECT 1261.880 2010.460 1262.140 2010.720 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 1261.880 3250.070 1262.140 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 1261.940 2010.750 1262.080 3250.070 ;
        RECT 1255.900 2010.430 1256.160 2010.750 ;
        RECT 1261.880 2010.430 1262.140 2010.750 ;
        RECT 1255.960 2000.000 1256.100 2010.430 ;
        RECT 1255.800 1999.540 1256.100 2000.000 ;
        RECT 1255.800 1996.000 1256.080 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1268.750 3484.900 1269.070 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 1268.750 3484.760 2901.150 3484.900 ;
        RECT 1268.750 3484.700 1269.070 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
        RECT 1263.690 2010.660 1264.010 2010.720 ;
        RECT 1268.750 2010.660 1269.070 2010.720 ;
        RECT 1263.690 2010.520 1269.070 2010.660 ;
        RECT 1263.690 2010.460 1264.010 2010.520 ;
        RECT 1268.750 2010.460 1269.070 2010.520 ;
      LAYER via ;
        RECT 1268.780 3484.700 1269.040 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
        RECT 1263.720 2010.460 1263.980 2010.720 ;
        RECT 1268.780 2010.460 1269.040 2010.720 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 1268.780 3484.670 1269.040 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 1268.840 2010.750 1268.980 3484.670 ;
        RECT 1263.720 2010.430 1263.980 2010.750 ;
        RECT 1268.780 2010.430 1269.040 2010.750 ;
        RECT 1263.780 2000.000 1263.920 2010.430 ;
        RECT 1263.620 1999.540 1263.920 2000.000 ;
        RECT 1263.620 1996.000 1263.900 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1276.110 3502.240 1276.430 3502.300 ;
        RECT 2635.870 3502.240 2636.190 3502.300 ;
        RECT 1276.110 3502.100 2636.190 3502.240 ;
        RECT 1276.110 3502.040 1276.430 3502.100 ;
        RECT 2635.870 3502.040 2636.190 3502.100 ;
        RECT 1271.970 2010.660 1272.290 2010.720 ;
        RECT 1276.110 2010.660 1276.430 2010.720 ;
        RECT 1271.970 2010.520 1276.430 2010.660 ;
        RECT 1271.970 2010.460 1272.290 2010.520 ;
        RECT 1276.110 2010.460 1276.430 2010.520 ;
      LAYER via ;
        RECT 1276.140 3502.040 1276.400 3502.300 ;
        RECT 2635.900 3502.040 2636.160 3502.300 ;
        RECT 1272.000 2010.460 1272.260 2010.720 ;
        RECT 1276.140 2010.460 1276.400 2010.720 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3502.330 2636.100 3517.600 ;
        RECT 1276.140 3502.010 1276.400 3502.330 ;
        RECT 2635.900 3502.010 2636.160 3502.330 ;
        RECT 1276.200 2010.750 1276.340 3502.010 ;
        RECT 1272.000 2010.430 1272.260 2010.750 ;
        RECT 1276.140 2010.430 1276.400 2010.750 ;
        RECT 1272.060 2000.000 1272.200 2010.430 ;
        RECT 1271.900 1999.540 1272.200 2000.000 ;
        RECT 1271.900 1996.000 1272.180 1999.540 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1282.090 3503.600 1282.410 3503.660 ;
        RECT 2311.570 3503.600 2311.890 3503.660 ;
        RECT 1282.090 3503.460 2311.890 3503.600 ;
        RECT 1282.090 3503.400 1282.410 3503.460 ;
        RECT 2311.570 3503.400 2311.890 3503.460 ;
      LAYER via ;
        RECT 1282.120 3503.400 1282.380 3503.660 ;
        RECT 2311.600 3503.400 2311.860 3503.660 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3503.690 2311.800 3517.600 ;
        RECT 1282.120 3503.370 1282.380 3503.690 ;
        RECT 2311.600 3503.370 2311.860 3503.690 ;
        RECT 1282.180 2001.650 1282.320 3503.370 ;
        RECT 1280.800 2001.510 1282.320 2001.650 ;
        RECT 1279.720 1999.610 1280.000 2000.000 ;
        RECT 1280.800 1999.610 1280.940 2001.510 ;
        RECT 1279.720 1999.470 1280.940 1999.610 ;
        RECT 1279.720 1996.000 1280.000 1999.470 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1289.450 3504.960 1289.770 3505.020 ;
        RECT 1987.270 3504.960 1987.590 3505.020 ;
        RECT 1289.450 3504.820 1987.590 3504.960 ;
        RECT 1289.450 3504.760 1289.770 3504.820 ;
        RECT 1987.270 3504.760 1987.590 3504.820 ;
      LAYER via ;
        RECT 1289.480 3504.760 1289.740 3505.020 ;
        RECT 1987.300 3504.760 1987.560 3505.020 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3505.050 1987.500 3517.600 ;
        RECT 1289.480 3504.730 1289.740 3505.050 ;
        RECT 1987.300 3504.730 1987.560 3505.050 ;
        RECT 1287.540 1999.610 1287.820 2000.000 ;
        RECT 1289.540 1999.610 1289.680 3504.730 ;
        RECT 1287.540 1999.470 1289.680 1999.610 ;
        RECT 1287.540 1996.000 1287.820 1999.470 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1295.890 3500.200 1296.210 3500.260 ;
        RECT 1662.510 3500.200 1662.830 3500.260 ;
        RECT 1295.890 3500.060 1662.830 3500.200 ;
        RECT 1295.890 3500.000 1296.210 3500.060 ;
        RECT 1662.510 3500.000 1662.830 3500.060 ;
      LAYER via ;
        RECT 1295.920 3500.000 1296.180 3500.260 ;
        RECT 1662.540 3500.000 1662.800 3500.260 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3500.290 1662.740 3517.600 ;
        RECT 1295.920 3499.970 1296.180 3500.290 ;
        RECT 1662.540 3499.970 1662.800 3500.290 ;
        RECT 1295.360 1999.610 1295.640 2000.000 ;
        RECT 1295.980 1999.610 1296.120 3499.970 ;
        RECT 1295.360 1999.470 1296.120 1999.610 ;
        RECT 1295.360 1996.000 1295.640 1999.470 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1303.710 3498.500 1304.030 3498.560 ;
        RECT 1338.210 3498.500 1338.530 3498.560 ;
        RECT 1303.710 3498.360 1338.530 3498.500 ;
        RECT 1303.710 3498.300 1304.030 3498.360 ;
        RECT 1338.210 3498.300 1338.530 3498.360 ;
      LAYER via ;
        RECT 1303.740 3498.300 1304.000 3498.560 ;
        RECT 1338.240 3498.300 1338.500 3498.560 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3498.590 1338.440 3517.600 ;
        RECT 1303.740 3498.270 1304.000 3498.590 ;
        RECT 1338.240 3498.270 1338.500 3498.590 ;
        RECT 1303.180 1999.610 1303.460 2000.000 ;
        RECT 1303.800 1999.610 1303.940 3498.270 ;
        RECT 1303.180 1999.470 1303.940 1999.610 ;
        RECT 1303.180 1996.000 1303.460 1999.470 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1177.285 1996.225 1177.455 1997.415 ;
      LAYER mcon ;
        RECT 1177.285 1997.245 1177.455 1997.415 ;
      LAYER met1 ;
        RECT 1162.490 1997.400 1162.810 1997.460 ;
        RECT 1177.225 1997.400 1177.515 1997.445 ;
        RECT 1162.490 1997.260 1177.515 1997.400 ;
        RECT 1162.490 1997.200 1162.810 1997.260 ;
        RECT 1177.225 1997.215 1177.515 1997.260 ;
        RECT 1177.225 1996.380 1177.515 1996.425 ;
        RECT 1528.190 1996.380 1528.510 1996.440 ;
        RECT 1177.225 1996.240 1528.510 1996.380 ;
        RECT 1177.225 1996.195 1177.515 1996.240 ;
        RECT 1528.190 1996.180 1528.510 1996.240 ;
        RECT 1528.190 441.560 1528.510 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 1528.190 441.420 2901.150 441.560 ;
        RECT 1528.190 441.360 1528.510 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 1162.520 1997.200 1162.780 1997.460 ;
        RECT 1528.220 1996.180 1528.480 1996.440 ;
        RECT 1528.220 441.360 1528.480 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 1161.040 1997.570 1161.320 2000.000 ;
        RECT 1161.040 1997.490 1162.720 1997.570 ;
        RECT 1161.040 1997.430 1162.780 1997.490 ;
        RECT 1161.040 1996.000 1161.320 1997.430 ;
        RECT 1162.520 1997.170 1162.780 1997.430 ;
        RECT 1528.220 1996.150 1528.480 1996.470 ;
        RECT 1528.280 441.650 1528.420 1996.150 ;
        RECT 1528.220 441.330 1528.480 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3499.860 1014.230 3499.920 ;
        RECT 1311.070 3499.860 1311.390 3499.920 ;
        RECT 1013.910 3499.720 1311.390 3499.860 ;
        RECT 1013.910 3499.660 1014.230 3499.720 ;
        RECT 1311.070 3499.660 1311.390 3499.720 ;
      LAYER via ;
        RECT 1013.940 3499.660 1014.200 3499.920 ;
        RECT 1311.100 3499.660 1311.360 3499.920 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3499.950 1014.140 3517.600 ;
        RECT 1013.940 3499.630 1014.200 3499.950 ;
        RECT 1311.100 3499.630 1311.360 3499.950 ;
        RECT 1311.160 2000.000 1311.300 3499.630 ;
        RECT 1311.000 1999.540 1311.300 2000.000 ;
        RECT 1311.000 1996.000 1311.280 1999.540 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.150 3501.220 689.470 3501.280 ;
        RECT 1318.890 3501.220 1319.210 3501.280 ;
        RECT 689.150 3501.080 1319.210 3501.220 ;
        RECT 689.150 3501.020 689.470 3501.080 ;
        RECT 1318.890 3501.020 1319.210 3501.080 ;
      LAYER via ;
        RECT 689.180 3501.020 689.440 3501.280 ;
        RECT 1318.920 3501.020 1319.180 3501.280 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3501.310 689.380 3517.600 ;
        RECT 689.180 3500.990 689.440 3501.310 ;
        RECT 1318.920 3500.990 1319.180 3501.310 ;
        RECT 1318.980 1999.610 1319.120 3500.990 ;
        RECT 1319.280 1999.610 1319.560 2000.000 ;
        RECT 1318.980 1999.470 1319.560 1999.610 ;
        RECT 1319.280 1996.000 1319.560 1999.470 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 3503.940 365.170 3504.000 ;
        RECT 1325.330 3503.940 1325.650 3504.000 ;
        RECT 364.850 3503.800 1325.650 3503.940 ;
        RECT 364.850 3503.740 365.170 3503.800 ;
        RECT 1325.330 3503.740 1325.650 3503.800 ;
      LAYER via ;
        RECT 364.880 3503.740 365.140 3504.000 ;
        RECT 1325.360 3503.740 1325.620 3504.000 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3504.030 365.080 3517.600 ;
        RECT 364.880 3503.710 365.140 3504.030 ;
        RECT 1325.360 3503.710 1325.620 3504.030 ;
        RECT 1325.420 1999.610 1325.560 3503.710 ;
        RECT 1327.100 1999.610 1327.380 2000.000 ;
        RECT 1325.420 1999.470 1327.380 1999.610 ;
        RECT 1327.100 1996.000 1327.380 1999.470 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 40.550 3502.580 40.870 3502.640 ;
        RECT 1332.690 3502.580 1333.010 3502.640 ;
        RECT 40.550 3502.440 1333.010 3502.580 ;
        RECT 40.550 3502.380 40.870 3502.440 ;
        RECT 1332.690 3502.380 1333.010 3502.440 ;
      LAYER via ;
        RECT 40.580 3502.380 40.840 3502.640 ;
        RECT 1332.720 3502.380 1332.980 3502.640 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3502.670 40.780 3517.600 ;
        RECT 40.580 3502.350 40.840 3502.670 ;
        RECT 1332.720 3502.350 1332.980 3502.670 ;
        RECT 1332.780 1999.610 1332.920 3502.350 ;
        RECT 1334.920 1999.610 1335.200 2000.000 ;
        RECT 1332.780 1999.470 1335.200 1999.610 ;
        RECT 1334.920 1996.000 1335.200 1999.470 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 1339.130 3263.900 1339.450 3263.960 ;
        RECT 15.250 3263.760 1339.450 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 1339.130 3263.700 1339.450 3263.760 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 1339.160 3263.700 1339.420 3263.960 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 1339.160 3263.670 1339.420 3263.990 ;
        RECT 1339.220 2011.170 1339.360 3263.670 ;
        RECT 1339.220 2011.030 1340.740 2011.170 ;
        RECT 1340.600 1998.930 1340.740 2011.030 ;
        RECT 1342.740 1998.930 1343.020 2000.000 ;
        RECT 1340.600 1998.790 1343.020 1998.930 ;
        RECT 1342.740 1996.000 1343.020 1998.790 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2974.220 16.950 2974.280 ;
        RECT 1346.490 2974.220 1346.810 2974.280 ;
        RECT 16.630 2974.080 1346.810 2974.220 ;
        RECT 16.630 2974.020 16.950 2974.080 ;
        RECT 1346.490 2974.020 1346.810 2974.080 ;
      LAYER via ;
        RECT 16.660 2974.020 16.920 2974.280 ;
        RECT 1346.520 2974.020 1346.780 2974.280 ;
      LAYER met2 ;
        RECT 16.650 2979.915 16.930 2980.285 ;
        RECT 16.720 2974.310 16.860 2979.915 ;
        RECT 16.660 2973.990 16.920 2974.310 ;
        RECT 1346.520 2973.990 1346.780 2974.310 ;
        RECT 1346.580 2000.290 1346.720 2973.990 ;
        RECT 1346.580 2000.150 1349.480 2000.290 ;
        RECT 1349.340 1999.610 1349.480 2000.150 ;
        RECT 1350.560 1999.610 1350.840 2000.000 ;
        RECT 1349.340 1999.470 1350.840 1999.610 ;
        RECT 1350.560 1996.000 1350.840 1999.470 ;
      LAYER via2 ;
        RECT 16.650 2979.960 16.930 2980.240 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.625 2980.250 16.955 2980.265 ;
        RECT -4.800 2979.950 16.955 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.625 2979.935 16.955 2979.950 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 2691.340 16.490 2691.400 ;
        RECT 1353.850 2691.340 1354.170 2691.400 ;
        RECT 16.170 2691.200 1354.170 2691.340 ;
        RECT 16.170 2691.140 16.490 2691.200 ;
        RECT 1353.850 2691.140 1354.170 2691.200 ;
      LAYER via ;
        RECT 16.200 2691.140 16.460 2691.400 ;
        RECT 1353.880 2691.140 1354.140 2691.400 ;
      LAYER met2 ;
        RECT 16.190 2692.955 16.470 2693.325 ;
        RECT 16.260 2691.430 16.400 2692.955 ;
        RECT 16.200 2691.110 16.460 2691.430 ;
        RECT 1353.880 2691.110 1354.140 2691.430 ;
        RECT 1353.940 2012.530 1354.080 2691.110 ;
        RECT 1353.940 2012.390 1357.760 2012.530 ;
        RECT 1357.620 1999.610 1357.760 2012.390 ;
        RECT 1358.380 1999.610 1358.660 2000.000 ;
        RECT 1357.620 1999.470 1358.660 1999.610 ;
        RECT 1358.380 1996.000 1358.660 1999.470 ;
      LAYER via2 ;
        RECT 16.190 2693.000 16.470 2693.280 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 16.165 2693.290 16.495 2693.305 ;
        RECT -4.800 2692.990 16.495 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 16.165 2692.975 16.495 2692.990 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 2401.320 15.110 2401.380 ;
        RECT 1362.590 2401.320 1362.910 2401.380 ;
        RECT 14.790 2401.180 1362.910 2401.320 ;
        RECT 14.790 2401.120 15.110 2401.180 ;
        RECT 1362.590 2401.120 1362.910 2401.180 ;
        RECT 1362.590 2010.320 1362.910 2010.380 ;
        RECT 1366.270 2010.320 1366.590 2010.380 ;
        RECT 1362.590 2010.180 1366.590 2010.320 ;
        RECT 1362.590 2010.120 1362.910 2010.180 ;
        RECT 1366.270 2010.120 1366.590 2010.180 ;
      LAYER via ;
        RECT 14.820 2401.120 15.080 2401.380 ;
        RECT 1362.620 2401.120 1362.880 2401.380 ;
        RECT 1362.620 2010.120 1362.880 2010.380 ;
        RECT 1366.300 2010.120 1366.560 2010.380 ;
      LAYER met2 ;
        RECT 14.810 2405.315 15.090 2405.685 ;
        RECT 14.880 2401.410 15.020 2405.315 ;
        RECT 14.820 2401.090 15.080 2401.410 ;
        RECT 1362.620 2401.090 1362.880 2401.410 ;
        RECT 1362.680 2010.410 1362.820 2401.090 ;
        RECT 1362.620 2010.090 1362.880 2010.410 ;
        RECT 1366.300 2010.090 1366.560 2010.410 ;
        RECT 1366.360 2000.000 1366.500 2010.090 ;
        RECT 1366.200 1999.540 1366.500 2000.000 ;
        RECT 1366.200 1996.000 1366.480 1999.540 ;
      LAYER via2 ;
        RECT 14.810 2405.360 15.090 2405.640 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 14.785 2405.650 15.115 2405.665 ;
        RECT -4.800 2405.350 15.115 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 14.785 2405.335 15.115 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2118.440 16.950 2118.500 ;
        RECT 1369.490 2118.440 1369.810 2118.500 ;
        RECT 16.630 2118.300 1369.810 2118.440 ;
        RECT 16.630 2118.240 16.950 2118.300 ;
        RECT 1369.490 2118.240 1369.810 2118.300 ;
        RECT 1369.490 2010.320 1369.810 2010.380 ;
        RECT 1374.550 2010.320 1374.870 2010.380 ;
        RECT 1369.490 2010.180 1374.870 2010.320 ;
        RECT 1369.490 2010.120 1369.810 2010.180 ;
        RECT 1374.550 2010.120 1374.870 2010.180 ;
      LAYER via ;
        RECT 16.660 2118.240 16.920 2118.500 ;
        RECT 1369.520 2118.240 1369.780 2118.500 ;
        RECT 1369.520 2010.120 1369.780 2010.380 ;
        RECT 1374.580 2010.120 1374.840 2010.380 ;
      LAYER met2 ;
        RECT 16.650 2118.355 16.930 2118.725 ;
        RECT 16.660 2118.210 16.920 2118.355 ;
        RECT 1369.520 2118.210 1369.780 2118.530 ;
        RECT 1369.580 2010.410 1369.720 2118.210 ;
        RECT 1369.520 2010.090 1369.780 2010.410 ;
        RECT 1374.580 2010.090 1374.840 2010.410 ;
        RECT 1374.640 2000.000 1374.780 2010.090 ;
        RECT 1374.480 1999.540 1374.780 2000.000 ;
        RECT 1374.480 1996.000 1374.760 1999.540 ;
      LAYER via2 ;
        RECT 16.650 2118.400 16.930 2118.680 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.625 2118.690 16.955 2118.705 ;
        RECT -4.800 2118.390 16.955 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.625 2118.375 16.955 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1134.890 2006.240 1135.210 2006.300 ;
        RECT 1382.370 2006.240 1382.690 2006.300 ;
        RECT 1134.890 2006.100 1382.690 2006.240 ;
        RECT 1134.890 2006.040 1135.210 2006.100 ;
        RECT 1382.370 2006.040 1382.690 2006.100 ;
        RECT 14.790 1835.220 15.110 1835.280 ;
        RECT 1134.890 1835.220 1135.210 1835.280 ;
        RECT 14.790 1835.080 1135.210 1835.220 ;
        RECT 14.790 1835.020 15.110 1835.080 ;
        RECT 1134.890 1835.020 1135.210 1835.080 ;
      LAYER via ;
        RECT 1134.920 2006.040 1135.180 2006.300 ;
        RECT 1382.400 2006.040 1382.660 2006.300 ;
        RECT 14.820 1835.020 15.080 1835.280 ;
        RECT 1134.920 1835.020 1135.180 1835.280 ;
      LAYER met2 ;
        RECT 1134.920 2006.010 1135.180 2006.330 ;
        RECT 1382.400 2006.010 1382.660 2006.330 ;
        RECT 1134.980 1835.310 1135.120 2006.010 ;
        RECT 1382.460 2000.000 1382.600 2006.010 ;
        RECT 1382.300 1999.540 1382.600 2000.000 ;
        RECT 1382.300 1996.000 1382.580 1999.540 ;
        RECT 14.820 1834.990 15.080 1835.310 ;
        RECT 1134.920 1834.990 1135.180 1835.310 ;
        RECT 14.880 1831.085 15.020 1834.990 ;
        RECT 14.810 1830.715 15.090 1831.085 ;
      LAYER via2 ;
        RECT 14.810 1830.760 15.090 1831.040 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 14.785 1831.050 15.115 1831.065 ;
        RECT -4.800 1830.750 15.115 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 14.785 1830.735 15.115 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1170.845 1994.865 1171.015 1996.395 ;
      LAYER mcon ;
        RECT 1170.845 1996.225 1171.015 1996.395 ;
      LAYER met1 ;
        RECT 1170.770 1996.380 1171.090 1996.440 ;
        RECT 1170.575 1996.240 1171.090 1996.380 ;
        RECT 1170.770 1996.180 1171.090 1996.240 ;
        RECT 1170.785 1995.020 1171.075 1995.065 ;
        RECT 1597.190 1995.020 1597.510 1995.080 ;
        RECT 1170.785 1994.880 1597.510 1995.020 ;
        RECT 1170.785 1994.835 1171.075 1994.880 ;
        RECT 1597.190 1994.820 1597.510 1994.880 ;
        RECT 1597.190 676.160 1597.510 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 1597.190 676.020 2901.150 676.160 ;
        RECT 1597.190 675.960 1597.510 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 1170.800 1996.180 1171.060 1996.440 ;
        RECT 1597.220 1994.820 1597.480 1995.080 ;
        RECT 1597.220 675.960 1597.480 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 1169.320 1996.890 1169.600 2000.000 ;
        RECT 1169.320 1996.750 1171.000 1996.890 ;
        RECT 1169.320 1996.000 1169.600 1996.750 ;
        RECT 1170.860 1996.470 1171.000 1996.750 ;
        RECT 1170.800 1996.150 1171.060 1996.470 ;
        RECT 1597.220 1994.790 1597.480 1995.110 ;
        RECT 1597.280 676.250 1597.420 1994.790 ;
        RECT 1597.220 675.930 1597.480 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1058.990 2003.520 1059.310 2003.580 ;
        RECT 1390.190 2003.520 1390.510 2003.580 ;
        RECT 1058.990 2003.380 1390.510 2003.520 ;
        RECT 1058.990 2003.320 1059.310 2003.380 ;
        RECT 1390.190 2003.320 1390.510 2003.380 ;
        RECT 17.090 1545.540 17.410 1545.600 ;
        RECT 1058.990 1545.540 1059.310 1545.600 ;
        RECT 17.090 1545.400 1059.310 1545.540 ;
        RECT 17.090 1545.340 17.410 1545.400 ;
        RECT 1058.990 1545.340 1059.310 1545.400 ;
      LAYER via ;
        RECT 1059.020 2003.320 1059.280 2003.580 ;
        RECT 1390.220 2003.320 1390.480 2003.580 ;
        RECT 17.120 1545.340 17.380 1545.600 ;
        RECT 1059.020 1545.340 1059.280 1545.600 ;
      LAYER met2 ;
        RECT 1059.020 2003.290 1059.280 2003.610 ;
        RECT 1390.220 2003.290 1390.480 2003.610 ;
        RECT 1059.080 1545.630 1059.220 2003.290 ;
        RECT 1390.280 2000.000 1390.420 2003.290 ;
        RECT 1390.120 1999.540 1390.420 2000.000 ;
        RECT 1390.120 1996.000 1390.400 1999.540 ;
        RECT 17.120 1545.310 17.380 1545.630 ;
        RECT 1059.020 1545.310 1059.280 1545.630 ;
        RECT 17.180 1544.125 17.320 1545.310 ;
        RECT 17.110 1543.755 17.390 1544.125 ;
      LAYER via2 ;
        RECT 17.110 1543.800 17.390 1544.080 ;
      LAYER met3 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 17.085 1544.090 17.415 1544.105 ;
        RECT -4.800 1543.790 17.415 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 17.085 1543.775 17.415 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1045.190 1996.720 1045.510 1996.780 ;
        RECT 1396.630 1996.720 1396.950 1996.780 ;
        RECT 1045.190 1996.580 1396.950 1996.720 ;
        RECT 1045.190 1996.520 1045.510 1996.580 ;
        RECT 1396.630 1996.520 1396.950 1996.580 ;
        RECT 14.330 1331.680 14.650 1331.740 ;
        RECT 1045.190 1331.680 1045.510 1331.740 ;
        RECT 14.330 1331.540 1045.510 1331.680 ;
        RECT 14.330 1331.480 14.650 1331.540 ;
        RECT 1045.190 1331.480 1045.510 1331.540 ;
      LAYER via ;
        RECT 1045.220 1996.520 1045.480 1996.780 ;
        RECT 1396.660 1996.520 1396.920 1996.780 ;
        RECT 14.360 1331.480 14.620 1331.740 ;
        RECT 1045.220 1331.480 1045.480 1331.740 ;
      LAYER met2 ;
        RECT 1397.940 1996.890 1398.220 2000.000 ;
        RECT 1396.720 1996.810 1398.220 1996.890 ;
        RECT 1045.220 1996.490 1045.480 1996.810 ;
        RECT 1396.660 1996.750 1398.220 1996.810 ;
        RECT 1396.660 1996.490 1396.920 1996.750 ;
        RECT 1045.280 1331.770 1045.420 1996.490 ;
        RECT 1397.940 1996.000 1398.220 1996.750 ;
        RECT 14.360 1331.450 14.620 1331.770 ;
        RECT 1045.220 1331.450 1045.480 1331.770 ;
        RECT 14.420 1328.565 14.560 1331.450 ;
        RECT 14.350 1328.195 14.630 1328.565 ;
      LAYER via2 ;
        RECT 14.350 1328.240 14.630 1328.520 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 14.325 1328.530 14.655 1328.545 ;
        RECT -4.800 1328.230 14.655 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 14.325 1328.215 14.655 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1038.290 2002.840 1038.610 2002.900 ;
        RECT 1405.830 2002.840 1406.150 2002.900 ;
        RECT 1038.290 2002.700 1406.150 2002.840 ;
        RECT 1038.290 2002.640 1038.610 2002.700 ;
        RECT 1405.830 2002.640 1406.150 2002.700 ;
        RECT 15.710 1117.820 16.030 1117.880 ;
        RECT 1038.290 1117.820 1038.610 1117.880 ;
        RECT 15.710 1117.680 1038.610 1117.820 ;
        RECT 15.710 1117.620 16.030 1117.680 ;
        RECT 1038.290 1117.620 1038.610 1117.680 ;
      LAYER via ;
        RECT 1038.320 2002.640 1038.580 2002.900 ;
        RECT 1405.860 2002.640 1406.120 2002.900 ;
        RECT 15.740 1117.620 16.000 1117.880 ;
        RECT 1038.320 1117.620 1038.580 1117.880 ;
      LAYER met2 ;
        RECT 1038.320 2002.610 1038.580 2002.930 ;
        RECT 1405.860 2002.610 1406.120 2002.930 ;
        RECT 1038.380 1117.910 1038.520 2002.610 ;
        RECT 1405.920 2000.000 1406.060 2002.610 ;
        RECT 1405.760 1999.540 1406.060 2000.000 ;
        RECT 1405.760 1996.000 1406.040 1999.540 ;
        RECT 15.740 1117.590 16.000 1117.910 ;
        RECT 1038.320 1117.590 1038.580 1117.910 ;
        RECT 15.800 1113.005 15.940 1117.590 ;
        RECT 15.730 1112.635 16.010 1113.005 ;
      LAYER via2 ;
        RECT 15.730 1112.680 16.010 1112.960 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 15.705 1112.970 16.035 1112.985 ;
        RECT -4.800 1112.670 16.035 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 15.705 1112.655 16.035 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1412.345 1995.545 1412.515 1996.735 ;
      LAYER mcon ;
        RECT 1412.345 1996.565 1412.515 1996.735 ;
      LAYER met1 ;
        RECT 1412.270 1996.720 1412.590 1996.780 ;
        RECT 1412.075 1996.580 1412.590 1996.720 ;
        RECT 1412.270 1996.520 1412.590 1996.580 ;
        RECT 1024.490 1995.700 1024.810 1995.760 ;
        RECT 1412.285 1995.700 1412.575 1995.745 ;
        RECT 1024.490 1995.560 1412.575 1995.700 ;
        RECT 1024.490 1995.500 1024.810 1995.560 ;
        RECT 1412.285 1995.515 1412.575 1995.560 ;
        RECT 16.170 903.960 16.490 904.020 ;
        RECT 1024.490 903.960 1024.810 904.020 ;
        RECT 16.170 903.820 1024.810 903.960 ;
        RECT 16.170 903.760 16.490 903.820 ;
        RECT 1024.490 903.760 1024.810 903.820 ;
      LAYER via ;
        RECT 1412.300 1996.520 1412.560 1996.780 ;
        RECT 1024.520 1995.500 1024.780 1995.760 ;
        RECT 16.200 903.760 16.460 904.020 ;
        RECT 1024.520 903.760 1024.780 904.020 ;
      LAYER met2 ;
        RECT 1413.580 1996.890 1413.860 2000.000 ;
        RECT 1412.360 1996.810 1413.860 1996.890 ;
        RECT 1412.300 1996.750 1413.860 1996.810 ;
        RECT 1412.300 1996.490 1412.560 1996.750 ;
        RECT 1413.580 1996.000 1413.860 1996.750 ;
        RECT 1024.520 1995.470 1024.780 1995.790 ;
        RECT 1024.580 904.050 1024.720 1995.470 ;
        RECT 16.200 903.730 16.460 904.050 ;
        RECT 1024.520 903.730 1024.780 904.050 ;
        RECT 16.260 897.445 16.400 903.730 ;
        RECT 16.190 897.075 16.470 897.445 ;
      LAYER via2 ;
        RECT 16.190 897.120 16.470 897.400 ;
      LAYER met3 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 16.165 897.410 16.495 897.425 ;
        RECT -4.800 897.110 16.495 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 16.165 897.095 16.495 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 682.960 16.490 683.020 ;
        RECT 86.090 682.960 86.410 683.020 ;
        RECT 16.170 682.820 86.410 682.960 ;
        RECT 16.170 682.760 16.490 682.820 ;
        RECT 86.090 682.760 86.410 682.820 ;
      LAYER via ;
        RECT 16.200 682.760 16.460 683.020 ;
        RECT 86.120 682.760 86.380 683.020 ;
      LAYER met2 ;
        RECT 1421.860 1996.890 1422.140 2000.000 ;
        RECT 1422.410 1996.890 1422.690 1997.005 ;
        RECT 1421.860 1996.750 1422.690 1996.890 ;
        RECT 1421.860 1996.000 1422.140 1996.750 ;
        RECT 1422.410 1996.635 1422.690 1996.750 ;
        RECT 86.110 1989.835 86.390 1990.205 ;
        RECT 86.180 683.050 86.320 1989.835 ;
        RECT 16.200 682.730 16.460 683.050 ;
        RECT 86.120 682.730 86.380 683.050 ;
        RECT 16.260 681.885 16.400 682.730 ;
        RECT 16.190 681.515 16.470 681.885 ;
      LAYER via2 ;
        RECT 1422.410 1996.680 1422.690 1996.960 ;
        RECT 86.110 1989.880 86.390 1990.160 ;
        RECT 16.190 681.560 16.470 681.840 ;
      LAYER met3 ;
        RECT 1421.670 1996.970 1422.050 1996.980 ;
        RECT 1422.385 1996.970 1422.715 1996.985 ;
        RECT 1421.670 1996.670 1422.715 1996.970 ;
        RECT 1421.670 1996.660 1422.050 1996.670 ;
        RECT 1422.385 1996.655 1422.715 1996.670 ;
        RECT 86.085 1990.170 86.415 1990.185 ;
        RECT 1421.670 1990.170 1422.050 1990.180 ;
        RECT 86.085 1989.870 1422.050 1990.170 ;
        RECT 86.085 1989.855 86.415 1989.870 ;
        RECT 1421.670 1989.860 1422.050 1989.870 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 16.165 681.850 16.495 681.865 ;
        RECT -4.800 681.550 16.495 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 16.165 681.535 16.495 681.550 ;
      LAYER via3 ;
        RECT 1421.700 1996.660 1422.020 1996.980 ;
        RECT 1421.700 1989.860 1422.020 1990.180 ;
      LAYER met4 ;
        RECT 1421.695 1996.655 1422.025 1996.985 ;
        RECT 1421.710 1990.185 1422.010 1996.655 ;
        RECT 1421.695 1989.855 1422.025 1990.185 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1017.590 2001.820 1017.910 2001.880 ;
        RECT 1429.750 2001.820 1430.070 2001.880 ;
        RECT 1017.590 2001.680 1430.070 2001.820 ;
        RECT 1017.590 2001.620 1017.910 2001.680 ;
        RECT 1429.750 2001.620 1430.070 2001.680 ;
        RECT 17.090 469.100 17.410 469.160 ;
        RECT 1017.590 469.100 1017.910 469.160 ;
        RECT 17.090 468.960 1017.910 469.100 ;
        RECT 17.090 468.900 17.410 468.960 ;
        RECT 1017.590 468.900 1017.910 468.960 ;
      LAYER via ;
        RECT 1017.620 2001.620 1017.880 2001.880 ;
        RECT 1429.780 2001.620 1430.040 2001.880 ;
        RECT 17.120 468.900 17.380 469.160 ;
        RECT 1017.620 468.900 1017.880 469.160 ;
      LAYER met2 ;
        RECT 1017.620 2001.590 1017.880 2001.910 ;
        RECT 1429.780 2001.590 1430.040 2001.910 ;
        RECT 1017.680 469.190 1017.820 2001.590 ;
        RECT 1429.840 2000.000 1429.980 2001.590 ;
        RECT 1429.680 1999.540 1429.980 2000.000 ;
        RECT 1429.680 1996.000 1429.960 1999.540 ;
        RECT 17.120 468.870 17.380 469.190 ;
        RECT 1017.620 468.870 1017.880 469.190 ;
        RECT 17.180 466.325 17.320 468.870 ;
        RECT 17.110 465.955 17.390 466.325 ;
      LAYER via2 ;
        RECT 17.110 466.000 17.390 466.280 ;
      LAYER met3 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.085 466.290 17.415 466.305 ;
        RECT -4.800 465.990 17.415 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.085 465.975 17.415 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 255.240 17.410 255.300 ;
        RECT 1003.790 255.240 1004.110 255.300 ;
        RECT 17.090 255.100 1004.110 255.240 ;
        RECT 17.090 255.040 17.410 255.100 ;
        RECT 1003.790 255.040 1004.110 255.100 ;
      LAYER via ;
        RECT 17.120 255.040 17.380 255.300 ;
        RECT 1003.820 255.040 1004.080 255.300 ;
      LAYER met2 ;
        RECT 1436.670 1996.890 1436.950 1997.005 ;
        RECT 1437.500 1996.890 1437.780 2000.000 ;
        RECT 1436.670 1996.750 1437.780 1996.890 ;
        RECT 1436.670 1996.635 1436.950 1996.750 ;
        RECT 1437.500 1996.000 1437.780 1996.750 ;
        RECT 1003.810 1991.195 1004.090 1991.565 ;
        RECT 1003.880 255.330 1004.020 1991.195 ;
        RECT 17.120 255.010 17.380 255.330 ;
        RECT 1003.820 255.010 1004.080 255.330 ;
        RECT 17.180 250.765 17.320 255.010 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 1436.670 1996.680 1436.950 1996.960 ;
        RECT 1003.810 1991.240 1004.090 1991.520 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
        RECT 1436.645 1996.980 1436.975 1996.985 ;
        RECT 1436.390 1996.970 1436.975 1996.980 ;
        RECT 1436.190 1996.670 1436.975 1996.970 ;
        RECT 1436.390 1996.660 1436.975 1996.670 ;
        RECT 1436.645 1996.655 1436.975 1996.660 ;
        RECT 1003.785 1991.530 1004.115 1991.545 ;
        RECT 1436.390 1991.530 1436.770 1991.540 ;
        RECT 1003.785 1991.230 1436.770 1991.530 ;
        RECT 1003.785 1991.215 1004.115 1991.230 ;
        RECT 1436.390 1991.220 1436.770 1991.230 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.085 250.415 17.415 250.430 ;
      LAYER via3 ;
        RECT 1436.420 1996.660 1436.740 1996.980 ;
        RECT 1436.420 1991.220 1436.740 1991.540 ;
      LAYER met4 ;
        RECT 1436.415 1996.655 1436.745 1996.985 ;
        RECT 1436.430 1991.545 1436.730 1996.655 ;
        RECT 1436.415 1991.215 1436.745 1991.545 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1443.625 1994.525 1443.795 1996.735 ;
      LAYER mcon ;
        RECT 1443.625 1996.565 1443.795 1996.735 ;
      LAYER met1 ;
        RECT 1443.550 1996.720 1443.870 1996.780 ;
        RECT 1443.355 1996.580 1443.870 1996.720 ;
        RECT 1443.550 1996.520 1443.870 1996.580 ;
        RECT 679.490 1994.680 679.810 1994.740 ;
        RECT 1443.565 1994.680 1443.855 1994.725 ;
        RECT 679.490 1994.540 1443.855 1994.680 ;
        RECT 679.490 1994.480 679.810 1994.540 ;
        RECT 1443.565 1994.495 1443.855 1994.540 ;
        RECT 17.090 41.380 17.410 41.440 ;
        RECT 679.490 41.380 679.810 41.440 ;
        RECT 17.090 41.240 679.810 41.380 ;
        RECT 17.090 41.180 17.410 41.240 ;
        RECT 679.490 41.180 679.810 41.240 ;
      LAYER via ;
        RECT 1443.580 1996.520 1443.840 1996.780 ;
        RECT 679.520 1994.480 679.780 1994.740 ;
        RECT 17.120 41.180 17.380 41.440 ;
        RECT 679.520 41.180 679.780 41.440 ;
      LAYER met2 ;
        RECT 1445.320 1996.890 1445.600 2000.000 ;
        RECT 1443.640 1996.810 1445.600 1996.890 ;
        RECT 1443.580 1996.750 1445.600 1996.810 ;
        RECT 1443.580 1996.490 1443.840 1996.750 ;
        RECT 1445.320 1996.000 1445.600 1996.750 ;
        RECT 679.520 1994.450 679.780 1994.770 ;
        RECT 679.580 41.470 679.720 1994.450 ;
        RECT 17.120 41.150 17.380 41.470 ;
        RECT 679.520 41.150 679.780 41.470 ;
        RECT 17.180 35.885 17.320 41.150 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1177.210 2002.160 1177.530 2002.220 ;
        RECT 1541.990 2002.160 1542.310 2002.220 ;
        RECT 1177.210 2002.020 1542.310 2002.160 ;
        RECT 1177.210 2001.960 1177.530 2002.020 ;
        RECT 1541.990 2001.960 1542.310 2002.020 ;
        RECT 1541.990 910.760 1542.310 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 1541.990 910.620 2901.150 910.760 ;
        RECT 1541.990 910.560 1542.310 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 1177.240 2001.960 1177.500 2002.220 ;
        RECT 1542.020 2001.960 1542.280 2002.220 ;
        RECT 1542.020 910.560 1542.280 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 1177.240 2001.930 1177.500 2002.250 ;
        RECT 1542.020 2001.930 1542.280 2002.250 ;
        RECT 1177.300 2000.000 1177.440 2001.930 ;
        RECT 1177.140 1999.540 1177.440 2000.000 ;
        RECT 1177.140 1996.000 1177.420 1999.540 ;
        RECT 1542.080 910.850 1542.220 2001.930 ;
        RECT 1542.020 910.530 1542.280 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2090.310 1139.920 2090.630 1139.980 ;
        RECT 2124.810 1139.920 2125.130 1139.980 ;
        RECT 2090.310 1139.780 2125.130 1139.920 ;
        RECT 2090.310 1139.720 2090.630 1139.780 ;
        RECT 2124.810 1139.720 2125.130 1139.780 ;
        RECT 2476.710 1139.580 2477.030 1139.640 ;
        RECT 2484.990 1139.580 2485.310 1139.640 ;
        RECT 2476.710 1139.440 2485.310 1139.580 ;
        RECT 2476.710 1139.380 2477.030 1139.440 ;
        RECT 2484.990 1139.380 2485.310 1139.440 ;
        RECT 2766.510 1139.580 2766.830 1139.640 ;
        RECT 2772.950 1139.580 2773.270 1139.640 ;
        RECT 2766.510 1139.440 2773.270 1139.580 ;
        RECT 2766.510 1139.380 2766.830 1139.440 ;
        RECT 2772.950 1139.380 2773.270 1139.440 ;
        RECT 2186.910 1139.240 2187.230 1139.300 ;
        RECT 2221.410 1139.240 2221.730 1139.300 ;
        RECT 2186.910 1139.100 2221.730 1139.240 ;
        RECT 2186.910 1139.040 2187.230 1139.100 ;
        RECT 2221.410 1139.040 2221.730 1139.100 ;
        RECT 2380.110 1139.240 2380.430 1139.300 ;
        RECT 2414.610 1139.240 2414.930 1139.300 ;
        RECT 2380.110 1139.100 2414.930 1139.240 ;
        RECT 2380.110 1139.040 2380.430 1139.100 ;
        RECT 2414.610 1139.040 2414.930 1139.100 ;
        RECT 2573.310 1139.240 2573.630 1139.300 ;
        RECT 2607.810 1139.240 2608.130 1139.300 ;
        RECT 2573.310 1139.100 2608.130 1139.240 ;
        RECT 2573.310 1139.040 2573.630 1139.100 ;
        RECT 2607.810 1139.040 2608.130 1139.100 ;
        RECT 1393.410 1138.900 1393.730 1138.960 ;
        RECT 1448.610 1138.900 1448.930 1138.960 ;
        RECT 1393.410 1138.760 1448.930 1138.900 ;
        RECT 1393.410 1138.700 1393.730 1138.760 ;
        RECT 1448.610 1138.700 1448.930 1138.760 ;
        RECT 1545.670 1138.900 1545.990 1138.960 ;
        RECT 1563.150 1138.900 1563.470 1138.960 ;
        RECT 1545.670 1138.760 1563.470 1138.900 ;
        RECT 1545.670 1138.700 1545.990 1138.760 ;
        RECT 1563.150 1138.700 1563.470 1138.760 ;
        RECT 2669.910 1138.900 2670.230 1138.960 ;
        RECT 2704.410 1138.900 2704.730 1138.960 ;
        RECT 2669.910 1138.760 2704.730 1138.900 ;
        RECT 2669.910 1138.700 2670.230 1138.760 ;
        RECT 2704.410 1138.700 2704.730 1138.760 ;
      LAYER via ;
        RECT 2090.340 1139.720 2090.600 1139.980 ;
        RECT 2124.840 1139.720 2125.100 1139.980 ;
        RECT 2476.740 1139.380 2477.000 1139.640 ;
        RECT 2485.020 1139.380 2485.280 1139.640 ;
        RECT 2766.540 1139.380 2766.800 1139.640 ;
        RECT 2772.980 1139.380 2773.240 1139.640 ;
        RECT 2186.940 1139.040 2187.200 1139.300 ;
        RECT 2221.440 1139.040 2221.700 1139.300 ;
        RECT 2380.140 1139.040 2380.400 1139.300 ;
        RECT 2414.640 1139.040 2414.900 1139.300 ;
        RECT 2573.340 1139.040 2573.600 1139.300 ;
        RECT 2607.840 1139.040 2608.100 1139.300 ;
        RECT 1393.440 1138.700 1393.700 1138.960 ;
        RECT 1448.640 1138.700 1448.900 1138.960 ;
        RECT 1545.700 1138.700 1545.960 1138.960 ;
        RECT 1563.180 1138.700 1563.440 1138.960 ;
        RECT 2669.940 1138.700 2670.200 1138.960 ;
        RECT 2704.440 1138.700 2704.700 1138.960 ;
      LAYER met2 ;
        RECT 1184.960 1996.890 1185.240 2000.000 ;
        RECT 1185.970 1996.890 1186.250 1997.005 ;
        RECT 1184.960 1996.750 1186.250 1996.890 ;
        RECT 1184.960 1996.000 1185.240 1996.750 ;
        RECT 1185.970 1996.635 1186.250 1996.750 ;
        RECT 1242.090 1139.835 1242.370 1140.205 ;
        RECT 1331.330 1139.835 1331.610 1140.205 ;
        RECT 1642.290 1140.090 1642.570 1140.205 ;
        RECT 1642.290 1139.950 1642.960 1140.090 ;
        RECT 1642.290 1139.835 1642.570 1139.950 ;
        RECT 1242.160 1139.525 1242.300 1139.835 ;
        RECT 1242.090 1139.155 1242.370 1139.525 ;
        RECT 1331.400 1138.845 1331.540 1139.835 ;
        RECT 1510.730 1139.155 1511.010 1139.525 ;
        RECT 1563.170 1139.155 1563.450 1139.525 ;
        RECT 1617.910 1139.155 1618.190 1139.525 ;
        RECT 1393.440 1138.845 1393.700 1138.990 ;
        RECT 1448.640 1138.845 1448.900 1138.990 ;
        RECT 1331.330 1138.475 1331.610 1138.845 ;
        RECT 1393.430 1138.475 1393.710 1138.845 ;
        RECT 1448.630 1138.475 1448.910 1138.845 ;
        RECT 1510.800 1137.485 1510.940 1139.155 ;
        RECT 1563.240 1138.990 1563.380 1139.155 ;
        RECT 1545.700 1138.845 1545.960 1138.990 ;
        RECT 1545.690 1138.475 1545.970 1138.845 ;
        RECT 1563.180 1138.670 1563.440 1138.990 ;
        RECT 1617.980 1138.165 1618.120 1139.155 ;
        RECT 1642.820 1138.165 1642.960 1139.950 ;
        RECT 2090.330 1139.835 2090.610 1140.205 ;
        RECT 2124.830 1139.835 2125.110 1140.205 ;
        RECT 2090.340 1139.690 2090.600 1139.835 ;
        RECT 2124.840 1139.690 2125.100 1139.835 ;
        RECT 2476.740 1139.525 2477.000 1139.670 ;
        RECT 2485.020 1139.525 2485.280 1139.670 ;
        RECT 2766.540 1139.525 2766.800 1139.670 ;
        RECT 2772.980 1139.525 2773.240 1139.670 ;
        RECT 2186.930 1139.155 2187.210 1139.525 ;
        RECT 2283.530 1139.410 2283.810 1139.525 ;
        RECT 2284.450 1139.410 2284.730 1139.525 ;
        RECT 2186.940 1139.010 2187.200 1139.155 ;
        RECT 2221.440 1139.010 2221.700 1139.330 ;
        RECT 2283.530 1139.270 2284.730 1139.410 ;
        RECT 2283.530 1139.155 2283.810 1139.270 ;
        RECT 2284.450 1139.155 2284.730 1139.270 ;
        RECT 2380.130 1139.155 2380.410 1139.525 ;
        RECT 2380.140 1139.010 2380.400 1139.155 ;
        RECT 2414.640 1139.010 2414.900 1139.330 ;
        RECT 2476.730 1139.155 2477.010 1139.525 ;
        RECT 2485.010 1139.155 2485.290 1139.525 ;
        RECT 2573.330 1139.155 2573.610 1139.525 ;
        RECT 2573.340 1139.010 2573.600 1139.155 ;
        RECT 2607.840 1139.010 2608.100 1139.330 ;
        RECT 2669.930 1139.155 2670.210 1139.525 ;
        RECT 2766.530 1139.155 2766.810 1139.525 ;
        RECT 2772.970 1139.155 2773.250 1139.525 ;
        RECT 2221.500 1138.845 2221.640 1139.010 ;
        RECT 2414.700 1138.845 2414.840 1139.010 ;
        RECT 2607.900 1138.845 2608.040 1139.010 ;
        RECT 2670.000 1138.990 2670.140 1139.155 ;
        RECT 2221.430 1138.475 2221.710 1138.845 ;
        RECT 2414.630 1138.475 2414.910 1138.845 ;
        RECT 2607.830 1138.475 2608.110 1138.845 ;
        RECT 2669.940 1138.670 2670.200 1138.990 ;
        RECT 2704.440 1138.845 2704.700 1138.990 ;
        RECT 2704.430 1138.475 2704.710 1138.845 ;
        RECT 1617.910 1137.795 1618.190 1138.165 ;
        RECT 1642.750 1137.795 1643.030 1138.165 ;
        RECT 1510.730 1137.115 1511.010 1137.485 ;
      LAYER via2 ;
        RECT 1185.970 1996.680 1186.250 1996.960 ;
        RECT 1242.090 1139.880 1242.370 1140.160 ;
        RECT 1331.330 1139.880 1331.610 1140.160 ;
        RECT 1642.290 1139.880 1642.570 1140.160 ;
        RECT 1242.090 1139.200 1242.370 1139.480 ;
        RECT 1510.730 1139.200 1511.010 1139.480 ;
        RECT 1563.170 1139.200 1563.450 1139.480 ;
        RECT 1617.910 1139.200 1618.190 1139.480 ;
        RECT 1331.330 1138.520 1331.610 1138.800 ;
        RECT 1393.430 1138.520 1393.710 1138.800 ;
        RECT 1448.630 1138.520 1448.910 1138.800 ;
        RECT 1545.690 1138.520 1545.970 1138.800 ;
        RECT 2090.330 1139.880 2090.610 1140.160 ;
        RECT 2124.830 1139.880 2125.110 1140.160 ;
        RECT 2186.930 1139.200 2187.210 1139.480 ;
        RECT 2283.530 1139.200 2283.810 1139.480 ;
        RECT 2284.450 1139.200 2284.730 1139.480 ;
        RECT 2380.130 1139.200 2380.410 1139.480 ;
        RECT 2476.730 1139.200 2477.010 1139.480 ;
        RECT 2485.010 1139.200 2485.290 1139.480 ;
        RECT 2573.330 1139.200 2573.610 1139.480 ;
        RECT 2669.930 1139.200 2670.210 1139.480 ;
        RECT 2766.530 1139.200 2766.810 1139.480 ;
        RECT 2772.970 1139.200 2773.250 1139.480 ;
        RECT 2221.430 1138.520 2221.710 1138.800 ;
        RECT 2414.630 1138.520 2414.910 1138.800 ;
        RECT 2607.830 1138.520 2608.110 1138.800 ;
        RECT 2704.430 1138.520 2704.710 1138.800 ;
        RECT 1617.910 1137.840 1618.190 1138.120 ;
        RECT 1642.750 1137.840 1643.030 1138.120 ;
        RECT 1510.730 1137.160 1511.010 1137.440 ;
      LAYER met3 ;
        RECT 1185.945 1996.980 1186.275 1996.985 ;
        RECT 1185.945 1996.970 1186.530 1996.980 ;
        RECT 1185.945 1996.670 1186.730 1996.970 ;
        RECT 1185.945 1996.660 1186.530 1996.670 ;
        RECT 1185.945 1996.655 1186.275 1996.660 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2916.710 1143.950 2924.800 1144.250 ;
        RECT 1242.065 1140.170 1242.395 1140.185 ;
        RECT 1331.305 1140.170 1331.635 1140.185 ;
        RECT 1642.265 1140.170 1642.595 1140.185 ;
        RECT 1242.065 1139.870 1331.635 1140.170 ;
        RECT 1242.065 1139.855 1242.395 1139.870 ;
        RECT 1331.305 1139.855 1331.635 1139.870 ;
        RECT 1641.590 1139.870 1642.595 1140.170 ;
        RECT 1186.150 1139.490 1186.530 1139.500 ;
        RECT 1242.065 1139.490 1242.395 1139.505 ;
        RECT 1510.705 1139.490 1511.035 1139.505 ;
        RECT 1186.150 1139.190 1242.395 1139.490 ;
        RECT 1186.150 1139.180 1186.530 1139.190 ;
        RECT 1242.065 1139.175 1242.395 1139.190 ;
        RECT 1463.110 1139.190 1511.035 1139.490 ;
        RECT 1331.305 1138.810 1331.635 1138.825 ;
        RECT 1393.405 1138.810 1393.735 1138.825 ;
        RECT 1331.305 1138.510 1393.735 1138.810 ;
        RECT 1331.305 1138.495 1331.635 1138.510 ;
        RECT 1393.405 1138.495 1393.735 1138.510 ;
        RECT 1448.605 1138.810 1448.935 1138.825 ;
        RECT 1463.110 1138.810 1463.410 1139.190 ;
        RECT 1510.705 1139.175 1511.035 1139.190 ;
        RECT 1563.145 1139.490 1563.475 1139.505 ;
        RECT 1593.710 1139.490 1594.090 1139.500 ;
        RECT 1563.145 1139.190 1594.090 1139.490 ;
        RECT 1563.145 1139.175 1563.475 1139.190 ;
        RECT 1593.710 1139.180 1594.090 1139.190 ;
        RECT 1617.885 1139.490 1618.215 1139.505 ;
        RECT 1641.590 1139.490 1641.890 1139.870 ;
        RECT 1642.265 1139.855 1642.595 1139.870 ;
        RECT 1690.310 1140.170 1690.690 1140.180 ;
        RECT 2090.305 1140.170 2090.635 1140.185 ;
        RECT 1690.310 1139.870 1773.450 1140.170 ;
        RECT 1690.310 1139.860 1690.690 1139.870 ;
        RECT 1617.885 1139.190 1641.890 1139.490 ;
        RECT 1773.150 1139.490 1773.450 1139.870 ;
        RECT 1821.910 1139.870 1870.050 1140.170 ;
        RECT 1773.150 1139.190 1821.290 1139.490 ;
        RECT 1617.885 1139.175 1618.215 1139.190 ;
        RECT 1545.665 1138.810 1545.995 1138.825 ;
        RECT 1690.310 1138.810 1690.690 1138.820 ;
        RECT 1448.605 1138.510 1463.410 1138.810 ;
        RECT 1544.990 1138.510 1545.995 1138.810 ;
        RECT 1448.605 1138.495 1448.935 1138.510 ;
        RECT 1510.705 1137.450 1511.035 1137.465 ;
        RECT 1544.990 1137.450 1545.290 1138.510 ;
        RECT 1545.665 1138.495 1545.995 1138.510 ;
        RECT 1657.230 1138.510 1690.690 1138.810 ;
        RECT 1820.990 1138.810 1821.290 1139.190 ;
        RECT 1821.910 1138.810 1822.210 1139.870 ;
        RECT 1869.750 1139.490 1870.050 1139.870 ;
        RECT 1918.510 1139.870 2041.170 1140.170 ;
        RECT 1869.750 1139.190 1917.890 1139.490 ;
        RECT 1820.990 1138.510 1822.210 1138.810 ;
        RECT 1917.590 1138.810 1917.890 1139.190 ;
        RECT 1918.510 1138.810 1918.810 1139.870 ;
        RECT 2040.870 1139.490 2041.170 1139.870 ;
        RECT 2076.750 1139.870 2090.635 1140.170 ;
        RECT 2076.750 1139.490 2077.050 1139.870 ;
        RECT 2090.305 1139.855 2090.635 1139.870 ;
        RECT 2124.805 1140.170 2125.135 1140.185 ;
        RECT 2124.805 1139.870 2138.690 1140.170 ;
        RECT 2124.805 1139.855 2125.135 1139.870 ;
        RECT 2040.870 1139.190 2077.050 1139.490 ;
        RECT 1917.590 1138.510 1918.810 1138.810 ;
        RECT 2138.390 1138.810 2138.690 1139.870 ;
        RECT 2186.905 1139.490 2187.235 1139.505 ;
        RECT 2283.505 1139.490 2283.835 1139.505 ;
        RECT 2139.310 1139.190 2187.235 1139.490 ;
        RECT 2139.310 1138.810 2139.610 1139.190 ;
        RECT 2186.905 1139.175 2187.235 1139.190 ;
        RECT 2235.910 1139.190 2283.835 1139.490 ;
        RECT 2138.390 1138.510 2139.610 1138.810 ;
        RECT 2221.405 1138.810 2221.735 1138.825 ;
        RECT 2235.910 1138.810 2236.210 1139.190 ;
        RECT 2283.505 1139.175 2283.835 1139.190 ;
        RECT 2284.425 1139.490 2284.755 1139.505 ;
        RECT 2380.105 1139.490 2380.435 1139.505 ;
        RECT 2476.705 1139.490 2477.035 1139.505 ;
        RECT 2284.425 1139.190 2331.890 1139.490 ;
        RECT 2284.425 1139.175 2284.755 1139.190 ;
        RECT 2221.405 1138.510 2236.210 1138.810 ;
        RECT 2331.590 1138.810 2331.890 1139.190 ;
        RECT 2332.510 1139.190 2380.435 1139.490 ;
        RECT 2332.510 1138.810 2332.810 1139.190 ;
        RECT 2380.105 1139.175 2380.435 1139.190 ;
        RECT 2429.110 1139.190 2477.035 1139.490 ;
        RECT 2331.590 1138.510 2332.810 1138.810 ;
        RECT 2414.605 1138.810 2414.935 1138.825 ;
        RECT 2429.110 1138.810 2429.410 1139.190 ;
        RECT 2476.705 1139.175 2477.035 1139.190 ;
        RECT 2484.985 1139.490 2485.315 1139.505 ;
        RECT 2573.305 1139.490 2573.635 1139.505 ;
        RECT 2669.905 1139.490 2670.235 1139.505 ;
        RECT 2766.505 1139.490 2766.835 1139.505 ;
        RECT 2484.985 1139.190 2525.090 1139.490 ;
        RECT 2484.985 1139.175 2485.315 1139.190 ;
        RECT 2414.605 1138.510 2429.410 1138.810 ;
        RECT 2524.790 1138.810 2525.090 1139.190 ;
        RECT 2525.710 1139.190 2573.635 1139.490 ;
        RECT 2525.710 1138.810 2526.010 1139.190 ;
        RECT 2573.305 1139.175 2573.635 1139.190 ;
        RECT 2622.310 1139.190 2670.235 1139.490 ;
        RECT 2524.790 1138.510 2526.010 1138.810 ;
        RECT 2607.805 1138.810 2608.135 1138.825 ;
        RECT 2622.310 1138.810 2622.610 1139.190 ;
        RECT 2669.905 1139.175 2670.235 1139.190 ;
        RECT 2718.910 1139.190 2766.835 1139.490 ;
        RECT 2607.805 1138.510 2622.610 1138.810 ;
        RECT 2704.405 1138.810 2704.735 1138.825 ;
        RECT 2718.910 1138.810 2719.210 1139.190 ;
        RECT 2766.505 1139.175 2766.835 1139.190 ;
        RECT 2772.945 1139.490 2773.275 1139.505 ;
        RECT 2916.710 1139.490 2917.010 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
        RECT 2772.945 1139.190 2814.890 1139.490 ;
        RECT 2772.945 1139.175 2773.275 1139.190 ;
        RECT 2704.405 1138.510 2719.210 1138.810 ;
        RECT 2814.590 1138.810 2814.890 1139.190 ;
        RECT 2884.510 1139.190 2917.010 1139.490 ;
        RECT 2884.510 1138.810 2884.810 1139.190 ;
        RECT 2814.590 1138.510 2884.810 1138.810 ;
        RECT 1593.710 1138.130 1594.090 1138.140 ;
        RECT 1617.885 1138.130 1618.215 1138.145 ;
        RECT 1593.710 1137.830 1618.215 1138.130 ;
        RECT 1593.710 1137.820 1594.090 1137.830 ;
        RECT 1617.885 1137.815 1618.215 1137.830 ;
        RECT 1642.725 1138.130 1643.055 1138.145 ;
        RECT 1657.230 1138.130 1657.530 1138.510 ;
        RECT 1690.310 1138.500 1690.690 1138.510 ;
        RECT 2221.405 1138.495 2221.735 1138.510 ;
        RECT 2414.605 1138.495 2414.935 1138.510 ;
        RECT 2607.805 1138.495 2608.135 1138.510 ;
        RECT 2704.405 1138.495 2704.735 1138.510 ;
        RECT 1642.725 1137.830 1657.530 1138.130 ;
        RECT 1642.725 1137.815 1643.055 1137.830 ;
        RECT 1510.705 1137.150 1545.290 1137.450 ;
        RECT 1510.705 1137.135 1511.035 1137.150 ;
      LAYER via3 ;
        RECT 1186.180 1996.660 1186.500 1996.980 ;
        RECT 1186.180 1139.180 1186.500 1139.500 ;
        RECT 1593.740 1139.180 1594.060 1139.500 ;
        RECT 1690.340 1139.860 1690.660 1140.180 ;
        RECT 1593.740 1137.820 1594.060 1138.140 ;
        RECT 1690.340 1138.500 1690.660 1138.820 ;
      LAYER met4 ;
        RECT 1186.175 1996.655 1186.505 1996.985 ;
        RECT 1186.190 1139.505 1186.490 1996.655 ;
        RECT 1690.335 1139.855 1690.665 1140.185 ;
        RECT 1186.175 1139.175 1186.505 1139.505 ;
        RECT 1593.735 1139.175 1594.065 1139.505 ;
        RECT 1593.750 1138.145 1594.050 1139.175 ;
        RECT 1690.350 1138.825 1690.650 1139.855 ;
        RECT 1690.335 1138.495 1690.665 1138.825 ;
        RECT 1593.735 1137.815 1594.065 1138.145 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1548.890 1379.960 1549.210 1380.020 ;
        RECT 2900.830 1379.960 2901.150 1380.020 ;
        RECT 1548.890 1379.820 2901.150 1379.960 ;
        RECT 1548.890 1379.760 1549.210 1379.820 ;
        RECT 2900.830 1379.760 2901.150 1379.820 ;
      LAYER via ;
        RECT 1548.920 1379.760 1549.180 1380.020 ;
        RECT 2900.860 1379.760 2901.120 1380.020 ;
      LAYER met2 ;
        RECT 1191.490 1996.890 1191.770 1997.005 ;
        RECT 1192.780 1996.890 1193.060 2000.000 ;
        RECT 1191.490 1996.750 1193.060 1996.890 ;
        RECT 1191.490 1996.635 1191.770 1996.750 ;
        RECT 1192.780 1996.000 1193.060 1996.750 ;
        RECT 1548.910 1992.555 1549.190 1992.925 ;
        RECT 1548.980 1380.050 1549.120 1992.555 ;
        RECT 1548.920 1379.730 1549.180 1380.050 ;
        RECT 2900.860 1379.730 2901.120 1380.050 ;
        RECT 2900.920 1378.885 2901.060 1379.730 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
      LAYER via2 ;
        RECT 1191.490 1996.680 1191.770 1996.960 ;
        RECT 1548.910 1992.600 1549.190 1992.880 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
      LAYER met3 ;
        RECT 1190.750 1996.970 1191.130 1996.980 ;
        RECT 1191.465 1996.970 1191.795 1996.985 ;
        RECT 1190.750 1996.670 1191.795 1996.970 ;
        RECT 1190.750 1996.660 1191.130 1996.670 ;
        RECT 1191.465 1996.655 1191.795 1996.670 ;
        RECT 1190.750 1992.890 1191.130 1992.900 ;
        RECT 1548.885 1992.890 1549.215 1992.905 ;
        RECT 1190.750 1992.590 1549.215 1992.890 ;
        RECT 1190.750 1992.580 1191.130 1992.590 ;
        RECT 1548.885 1992.575 1549.215 1992.590 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
      LAYER via3 ;
        RECT 1190.780 1996.660 1191.100 1996.980 ;
        RECT 1190.780 1992.580 1191.100 1992.900 ;
      LAYER met4 ;
        RECT 1190.775 1996.655 1191.105 1996.985 ;
        RECT 1190.790 1992.905 1191.090 1996.655 ;
        RECT 1190.775 1992.575 1191.105 1992.905 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1200.670 2001.140 1200.990 2001.200 ;
        RECT 1452.750 2001.140 1453.070 2001.200 ;
        RECT 1200.670 2001.000 1453.070 2001.140 ;
        RECT 1200.670 2000.940 1200.990 2001.000 ;
        RECT 1452.750 2000.940 1453.070 2001.000 ;
        RECT 1452.750 1614.560 1453.070 1614.620 ;
        RECT 2900.830 1614.560 2901.150 1614.620 ;
        RECT 1452.750 1614.420 2901.150 1614.560 ;
        RECT 1452.750 1614.360 1453.070 1614.420 ;
        RECT 2900.830 1614.360 2901.150 1614.420 ;
      LAYER via ;
        RECT 1200.700 2000.940 1200.960 2001.200 ;
        RECT 1452.780 2000.940 1453.040 2001.200 ;
        RECT 1452.780 1614.360 1453.040 1614.620 ;
        RECT 2900.860 1614.360 2901.120 1614.620 ;
      LAYER met2 ;
        RECT 1200.700 2000.910 1200.960 2001.230 ;
        RECT 1452.780 2000.910 1453.040 2001.230 ;
        RECT 1200.760 2000.000 1200.900 2000.910 ;
        RECT 1200.600 1999.540 1200.900 2000.000 ;
        RECT 1200.600 1996.000 1200.880 1999.540 ;
        RECT 1452.840 1614.650 1452.980 2000.910 ;
        RECT 1452.780 1614.330 1453.040 1614.650 ;
        RECT 2900.860 1614.330 2901.120 1614.650 ;
        RECT 2900.920 1613.485 2901.060 1614.330 ;
        RECT 2900.850 1613.115 2901.130 1613.485 ;
      LAYER via2 ;
        RECT 2900.850 1613.160 2901.130 1613.440 ;
      LAYER met3 ;
        RECT 2900.825 1613.450 2901.155 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2900.825 1613.150 2924.800 1613.450 ;
        RECT 2900.825 1613.135 2901.155 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1210.405 1994.185 1210.575 1999.455 ;
      LAYER mcon ;
        RECT 1210.405 1999.285 1210.575 1999.455 ;
      LAYER met1 ;
        RECT 1210.330 1999.440 1210.650 1999.500 ;
        RECT 1210.135 1999.300 1210.650 1999.440 ;
        RECT 1210.330 1999.240 1210.650 1999.300 ;
        RECT 1210.345 1994.340 1210.635 1994.385 ;
        RECT 1459.190 1994.340 1459.510 1994.400 ;
        RECT 1210.345 1994.200 1459.510 1994.340 ;
        RECT 1210.345 1994.155 1210.635 1994.200 ;
        RECT 1459.190 1994.140 1459.510 1994.200 ;
        RECT 1459.190 1849.160 1459.510 1849.220 ;
        RECT 2900.830 1849.160 2901.150 1849.220 ;
        RECT 1459.190 1849.020 2901.150 1849.160 ;
        RECT 1459.190 1848.960 1459.510 1849.020 ;
        RECT 2900.830 1848.960 2901.150 1849.020 ;
      LAYER via ;
        RECT 1210.360 1999.240 1210.620 1999.500 ;
        RECT 1459.220 1994.140 1459.480 1994.400 ;
        RECT 1459.220 1848.960 1459.480 1849.220 ;
        RECT 2900.860 1848.960 2901.120 1849.220 ;
      LAYER met2 ;
        RECT 1208.420 1999.610 1208.700 2000.000 ;
        RECT 1208.420 1999.530 1210.560 1999.610 ;
        RECT 1208.420 1999.470 1210.620 1999.530 ;
        RECT 1208.420 1996.000 1208.700 1999.470 ;
        RECT 1210.360 1999.210 1210.620 1999.470 ;
        RECT 1459.220 1994.110 1459.480 1994.430 ;
        RECT 1459.280 1849.250 1459.420 1994.110 ;
        RECT 1459.220 1848.930 1459.480 1849.250 ;
        RECT 2900.860 1848.930 2901.120 1849.250 ;
        RECT 2900.920 1848.085 2901.060 1848.930 ;
        RECT 2900.850 1847.715 2901.130 1848.085 ;
      LAYER via2 ;
        RECT 2900.850 1847.760 2901.130 1848.040 ;
      LAYER met3 ;
        RECT 2900.825 1848.050 2901.155 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2900.825 1847.750 2924.800 1848.050 ;
        RECT 2900.825 1847.735 2901.155 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1220.910 2077.300 1221.230 2077.360 ;
        RECT 2900.830 2077.300 2901.150 2077.360 ;
        RECT 1220.910 2077.160 2901.150 2077.300 ;
        RECT 1220.910 2077.100 1221.230 2077.160 ;
        RECT 2900.830 2077.100 2901.150 2077.160 ;
        RECT 1216.310 2009.300 1216.630 2009.360 ;
        RECT 1220.910 2009.300 1221.230 2009.360 ;
        RECT 1216.310 2009.160 1221.230 2009.300 ;
        RECT 1216.310 2009.100 1216.630 2009.160 ;
        RECT 1220.910 2009.100 1221.230 2009.160 ;
      LAYER via ;
        RECT 1220.940 2077.100 1221.200 2077.360 ;
        RECT 2900.860 2077.100 2901.120 2077.360 ;
        RECT 1216.340 2009.100 1216.600 2009.360 ;
        RECT 1220.940 2009.100 1221.200 2009.360 ;
      LAYER met2 ;
        RECT 2900.850 2082.315 2901.130 2082.685 ;
        RECT 2900.920 2077.390 2901.060 2082.315 ;
        RECT 1220.940 2077.070 1221.200 2077.390 ;
        RECT 2900.860 2077.070 2901.120 2077.390 ;
        RECT 1221.000 2009.390 1221.140 2077.070 ;
        RECT 1216.340 2009.070 1216.600 2009.390 ;
        RECT 1220.940 2009.070 1221.200 2009.390 ;
        RECT 1216.400 2000.000 1216.540 2009.070 ;
        RECT 1216.240 1999.540 1216.540 2000.000 ;
        RECT 1216.240 1996.000 1216.520 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2082.360 2901.130 2082.640 ;
      LAYER met3 ;
        RECT 2900.825 2082.650 2901.155 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.825 2082.350 2924.800 2082.650 ;
        RECT 2900.825 2082.335 2901.155 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 2311.900 1228.130 2311.960 ;
        RECT 2900.830 2311.900 2901.150 2311.960 ;
        RECT 1227.810 2311.760 2901.150 2311.900 ;
        RECT 1227.810 2311.700 1228.130 2311.760 ;
        RECT 2900.830 2311.700 2901.150 2311.760 ;
        RECT 1224.590 2009.640 1224.910 2009.700 ;
        RECT 1227.810 2009.640 1228.130 2009.700 ;
        RECT 1224.590 2009.500 1228.130 2009.640 ;
        RECT 1224.590 2009.440 1224.910 2009.500 ;
        RECT 1227.810 2009.440 1228.130 2009.500 ;
      LAYER via ;
        RECT 1227.840 2311.700 1228.100 2311.960 ;
        RECT 2900.860 2311.700 2901.120 2311.960 ;
        RECT 1224.620 2009.440 1224.880 2009.700 ;
        RECT 1227.840 2009.440 1228.100 2009.700 ;
      LAYER met2 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
        RECT 2900.920 2311.990 2901.060 2316.915 ;
        RECT 1227.840 2311.670 1228.100 2311.990 ;
        RECT 2900.860 2311.670 2901.120 2311.990 ;
        RECT 1227.900 2009.730 1228.040 2311.670 ;
        RECT 1224.620 2009.410 1224.880 2009.730 ;
        RECT 1227.840 2009.410 1228.100 2009.730 ;
        RECT 1224.680 2000.000 1224.820 2009.410 ;
        RECT 1224.520 1999.540 1224.820 2000.000 ;
        RECT 1224.520 1996.000 1224.800 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
      LAYER met3 ;
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1990.490 146.440 1990.810 146.500 ;
        RECT 2028.210 146.440 2028.530 146.500 ;
        RECT 1990.490 146.300 2028.530 146.440 ;
        RECT 1990.490 146.240 1990.810 146.300 ;
        RECT 2028.210 146.240 2028.530 146.300 ;
        RECT 2183.690 146.440 2184.010 146.500 ;
        RECT 2221.410 146.440 2221.730 146.500 ;
        RECT 2183.690 146.300 2221.730 146.440 ;
        RECT 2183.690 146.240 2184.010 146.300 ;
        RECT 2221.410 146.240 2221.730 146.300 ;
        RECT 2086.630 146.100 2086.950 146.160 ;
        RECT 2124.810 146.100 2125.130 146.160 ;
        RECT 2086.630 145.960 2125.130 146.100 ;
        RECT 2086.630 145.900 2086.950 145.960 ;
        RECT 2124.810 145.900 2125.130 145.960 ;
        RECT 2283.510 146.100 2283.830 146.160 ;
        RECT 2318.010 146.100 2318.330 146.160 ;
        RECT 2283.510 145.960 2318.330 146.100 ;
        RECT 2283.510 145.900 2283.830 145.960 ;
        RECT 2318.010 145.900 2318.330 145.960 ;
        RECT 2376.430 146.100 2376.750 146.160 ;
        RECT 2414.610 146.100 2414.930 146.160 ;
        RECT 2376.430 145.960 2414.930 146.100 ;
        RECT 2376.430 145.900 2376.750 145.960 ;
        RECT 2414.610 145.900 2414.930 145.960 ;
        RECT 2475.790 146.100 2476.110 146.160 ;
        RECT 2511.210 146.100 2511.530 146.160 ;
        RECT 2475.790 145.960 2511.530 146.100 ;
        RECT 2475.790 145.900 2476.110 145.960 ;
        RECT 2511.210 145.900 2511.530 145.960 ;
        RECT 2567.790 146.100 2568.110 146.160 ;
        RECT 2607.810 146.100 2608.130 146.160 ;
        RECT 2567.790 145.960 2608.130 146.100 ;
        RECT 2567.790 145.900 2568.110 145.960 ;
        RECT 2607.810 145.900 2608.130 145.960 ;
        RECT 2668.990 146.100 2669.310 146.160 ;
        RECT 2704.410 146.100 2704.730 146.160 ;
        RECT 2668.990 145.960 2704.730 146.100 ;
        RECT 2668.990 145.900 2669.310 145.960 ;
        RECT 2704.410 145.900 2704.730 145.960 ;
        RECT 2762.370 146.100 2762.690 146.160 ;
        RECT 2801.010 146.100 2801.330 146.160 ;
        RECT 2762.370 145.960 2801.330 146.100 ;
        RECT 2762.370 145.900 2762.690 145.960 ;
        RECT 2801.010 145.900 2801.330 145.960 ;
        RECT 1401.230 145.420 1401.550 145.480 ;
        RECT 1448.610 145.420 1448.930 145.480 ;
        RECT 1401.230 145.280 1448.930 145.420 ;
        RECT 1401.230 145.220 1401.550 145.280 ;
        RECT 1448.610 145.220 1448.930 145.280 ;
      LAYER via ;
        RECT 1990.520 146.240 1990.780 146.500 ;
        RECT 2028.240 146.240 2028.500 146.500 ;
        RECT 2183.720 146.240 2183.980 146.500 ;
        RECT 2221.440 146.240 2221.700 146.500 ;
        RECT 2086.660 145.900 2086.920 146.160 ;
        RECT 2124.840 145.900 2125.100 146.160 ;
        RECT 2283.540 145.900 2283.800 146.160 ;
        RECT 2318.040 145.900 2318.300 146.160 ;
        RECT 2376.460 145.900 2376.720 146.160 ;
        RECT 2414.640 145.900 2414.900 146.160 ;
        RECT 2475.820 145.900 2476.080 146.160 ;
        RECT 2511.240 145.900 2511.500 146.160 ;
        RECT 2567.820 145.900 2568.080 146.160 ;
        RECT 2607.840 145.900 2608.100 146.160 ;
        RECT 2669.020 145.900 2669.280 146.160 ;
        RECT 2704.440 145.900 2704.700 146.160 ;
        RECT 2762.400 145.900 2762.660 146.160 ;
        RECT 2801.040 145.900 2801.300 146.160 ;
        RECT 1401.260 145.220 1401.520 145.480 ;
        RECT 1448.640 145.220 1448.900 145.480 ;
      LAYER met2 ;
        RECT 1155.980 1996.890 1156.260 2000.000 ;
        RECT 1157.910 1996.890 1158.190 1997.005 ;
        RECT 1155.980 1996.750 1158.190 1996.890 ;
        RECT 1155.980 1996.000 1156.260 1996.750 ;
        RECT 1157.910 1996.635 1158.190 1996.750 ;
        RECT 1990.520 146.210 1990.780 146.530 ;
        RECT 2028.230 146.355 2028.510 146.725 ;
        RECT 2124.830 146.355 2125.110 146.725 ;
        RECT 2028.240 146.210 2028.500 146.355 ;
        RECT 1990.580 146.045 1990.720 146.210 ;
        RECT 2124.900 146.190 2125.040 146.355 ;
        RECT 2183.720 146.210 2183.980 146.530 ;
        RECT 2221.430 146.355 2221.710 146.725 ;
        RECT 2318.030 146.355 2318.310 146.725 ;
        RECT 2414.630 146.355 2414.910 146.725 ;
        RECT 2511.230 146.355 2511.510 146.725 ;
        RECT 2607.830 146.355 2608.110 146.725 ;
        RECT 2704.430 146.355 2704.710 146.725 ;
        RECT 2801.030 146.355 2801.310 146.725 ;
        RECT 2221.440 146.210 2221.700 146.355 ;
        RECT 2086.660 146.045 2086.920 146.190 ;
        RECT 1990.510 145.675 1990.790 146.045 ;
        RECT 2086.650 145.675 2086.930 146.045 ;
        RECT 2124.840 145.870 2125.100 146.190 ;
        RECT 2183.780 146.045 2183.920 146.210 ;
        RECT 2318.100 146.190 2318.240 146.355 ;
        RECT 2414.700 146.190 2414.840 146.355 ;
        RECT 2511.300 146.190 2511.440 146.355 ;
        RECT 2607.900 146.190 2608.040 146.355 ;
        RECT 2704.500 146.190 2704.640 146.355 ;
        RECT 2801.100 146.190 2801.240 146.355 ;
        RECT 2283.540 146.045 2283.800 146.190 ;
        RECT 2183.710 145.675 2183.990 146.045 ;
        RECT 2283.530 145.675 2283.810 146.045 ;
        RECT 2318.040 145.870 2318.300 146.190 ;
        RECT 2376.460 146.045 2376.720 146.190 ;
        RECT 2376.450 145.675 2376.730 146.045 ;
        RECT 2414.640 145.870 2414.900 146.190 ;
        RECT 2475.820 146.045 2476.080 146.190 ;
        RECT 2475.810 145.675 2476.090 146.045 ;
        RECT 2511.240 145.870 2511.500 146.190 ;
        RECT 2567.820 146.045 2568.080 146.190 ;
        RECT 2567.810 145.675 2568.090 146.045 ;
        RECT 2607.840 145.870 2608.100 146.190 ;
        RECT 2669.020 146.045 2669.280 146.190 ;
        RECT 2669.010 145.675 2669.290 146.045 ;
        RECT 2704.440 145.870 2704.700 146.190 ;
        RECT 2762.400 146.045 2762.660 146.190 ;
        RECT 2762.390 145.675 2762.670 146.045 ;
        RECT 2801.040 145.870 2801.300 146.190 ;
        RECT 1401.260 145.365 1401.520 145.510 ;
        RECT 1448.640 145.365 1448.900 145.510 ;
        RECT 1401.250 144.995 1401.530 145.365 ;
        RECT 1448.630 144.995 1448.910 145.365 ;
      LAYER via2 ;
        RECT 1157.910 1996.680 1158.190 1996.960 ;
        RECT 2028.230 146.400 2028.510 146.680 ;
        RECT 2124.830 146.400 2125.110 146.680 ;
        RECT 2221.430 146.400 2221.710 146.680 ;
        RECT 2318.030 146.400 2318.310 146.680 ;
        RECT 2414.630 146.400 2414.910 146.680 ;
        RECT 2511.230 146.400 2511.510 146.680 ;
        RECT 2607.830 146.400 2608.110 146.680 ;
        RECT 2704.430 146.400 2704.710 146.680 ;
        RECT 2801.030 146.400 2801.310 146.680 ;
        RECT 1990.510 145.720 1990.790 146.000 ;
        RECT 2086.650 145.720 2086.930 146.000 ;
        RECT 2183.710 145.720 2183.990 146.000 ;
        RECT 2283.530 145.720 2283.810 146.000 ;
        RECT 2376.450 145.720 2376.730 146.000 ;
        RECT 2475.810 145.720 2476.090 146.000 ;
        RECT 2567.810 145.720 2568.090 146.000 ;
        RECT 2669.010 145.720 2669.290 146.000 ;
        RECT 2762.390 145.720 2762.670 146.000 ;
        RECT 1401.250 145.040 1401.530 145.320 ;
        RECT 1448.630 145.040 1448.910 145.320 ;
      LAYER met3 ;
        RECT 1157.885 1996.970 1158.215 1996.985 ;
        RECT 1158.550 1996.970 1158.930 1996.980 ;
        RECT 1157.885 1996.670 1158.930 1996.970 ;
        RECT 1157.885 1996.655 1158.215 1996.670 ;
        RECT 1158.550 1996.660 1158.930 1996.670 ;
        RECT 1181.590 147.070 1255.490 147.370 ;
        RECT 1158.550 145.330 1158.930 145.340 ;
        RECT 1181.590 145.330 1181.890 147.070 ;
        RECT 1158.550 145.030 1181.890 145.330 ;
        RECT 1255.190 145.330 1255.490 147.070 ;
        RECT 2028.205 146.690 2028.535 146.705 ;
        RECT 2124.805 146.690 2125.135 146.705 ;
        RECT 2221.405 146.690 2221.735 146.705 ;
        RECT 2318.005 146.690 2318.335 146.705 ;
        RECT 2414.605 146.690 2414.935 146.705 ;
        RECT 2511.205 146.690 2511.535 146.705 ;
        RECT 2607.805 146.690 2608.135 146.705 ;
        RECT 2704.405 146.690 2704.735 146.705 ;
        RECT 2801.005 146.690 2801.335 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 1510.950 146.390 1607.850 146.690 ;
        RECT 1401.225 145.330 1401.555 145.345 ;
        RECT 1255.190 145.030 1401.555 145.330 ;
        RECT 1158.550 145.020 1158.930 145.030 ;
        RECT 1401.225 145.015 1401.555 145.030 ;
        RECT 1448.605 145.330 1448.935 145.345 ;
        RECT 1510.950 145.330 1511.250 146.390 ;
        RECT 1607.550 146.010 1607.850 146.390 ;
        RECT 1676.550 146.390 1724.690 146.690 ;
        RECT 1607.550 145.710 1655.690 146.010 ;
        RECT 1448.605 145.030 1511.250 145.330 ;
        RECT 1655.390 145.330 1655.690 145.710 ;
        RECT 1676.550 145.330 1676.850 146.390 ;
        RECT 1655.390 145.030 1676.850 145.330 ;
        RECT 1724.390 145.330 1724.690 146.390 ;
        RECT 1725.310 146.390 1773.450 146.690 ;
        RECT 1725.310 145.330 1725.610 146.390 ;
        RECT 1773.150 146.010 1773.450 146.390 ;
        RECT 1821.910 146.390 1870.050 146.690 ;
        RECT 1773.150 145.710 1821.290 146.010 ;
        RECT 1724.390 145.030 1725.610 145.330 ;
        RECT 1820.990 145.330 1821.290 145.710 ;
        RECT 1821.910 145.330 1822.210 146.390 ;
        RECT 1869.750 146.010 1870.050 146.390 ;
        RECT 1918.510 146.390 1946.410 146.690 ;
        RECT 1869.750 145.710 1917.890 146.010 ;
        RECT 1820.990 145.030 1822.210 145.330 ;
        RECT 1917.590 145.330 1917.890 145.710 ;
        RECT 1918.510 145.330 1918.810 146.390 ;
        RECT 1946.110 146.010 1946.410 146.390 ;
        RECT 2028.205 146.390 2043.010 146.690 ;
        RECT 2028.205 146.375 2028.535 146.390 ;
        RECT 1990.485 146.010 1990.815 146.025 ;
        RECT 1946.110 145.710 1990.815 146.010 ;
        RECT 2042.710 146.010 2043.010 146.390 ;
        RECT 2124.805 146.390 2139.610 146.690 ;
        RECT 2124.805 146.375 2125.135 146.390 ;
        RECT 2086.625 146.010 2086.955 146.025 ;
        RECT 2042.710 145.710 2086.955 146.010 ;
        RECT 2139.310 146.010 2139.610 146.390 ;
        RECT 2221.405 146.390 2236.210 146.690 ;
        RECT 2221.405 146.375 2221.735 146.390 ;
        RECT 2183.685 146.010 2184.015 146.025 ;
        RECT 2139.310 145.710 2184.015 146.010 ;
        RECT 2235.910 146.010 2236.210 146.390 ;
        RECT 2318.005 146.390 2332.810 146.690 ;
        RECT 2318.005 146.375 2318.335 146.390 ;
        RECT 2283.505 146.010 2283.835 146.025 ;
        RECT 2235.910 145.710 2283.835 146.010 ;
        RECT 2332.510 146.010 2332.810 146.390 ;
        RECT 2414.605 146.390 2429.410 146.690 ;
        RECT 2414.605 146.375 2414.935 146.390 ;
        RECT 2376.425 146.010 2376.755 146.025 ;
        RECT 2332.510 145.710 2376.755 146.010 ;
        RECT 2429.110 146.010 2429.410 146.390 ;
        RECT 2511.205 146.390 2526.010 146.690 ;
        RECT 2511.205 146.375 2511.535 146.390 ;
        RECT 2475.785 146.010 2476.115 146.025 ;
        RECT 2429.110 145.710 2476.115 146.010 ;
        RECT 2525.710 146.010 2526.010 146.390 ;
        RECT 2607.805 146.390 2622.610 146.690 ;
        RECT 2607.805 146.375 2608.135 146.390 ;
        RECT 2567.785 146.010 2568.115 146.025 ;
        RECT 2525.710 145.710 2568.115 146.010 ;
        RECT 2622.310 146.010 2622.610 146.390 ;
        RECT 2704.405 146.390 2719.210 146.690 ;
        RECT 2704.405 146.375 2704.735 146.390 ;
        RECT 2668.985 146.010 2669.315 146.025 ;
        RECT 2622.310 145.710 2669.315 146.010 ;
        RECT 2718.910 146.010 2719.210 146.390 ;
        RECT 2801.005 146.390 2863.650 146.690 ;
        RECT 2801.005 146.375 2801.335 146.390 ;
        RECT 2762.365 146.010 2762.695 146.025 ;
        RECT 2718.910 145.710 2762.695 146.010 ;
        RECT 1990.485 145.695 1990.815 145.710 ;
        RECT 2086.625 145.695 2086.955 145.710 ;
        RECT 2183.685 145.695 2184.015 145.710 ;
        RECT 2283.505 145.695 2283.835 145.710 ;
        RECT 2376.425 145.695 2376.755 145.710 ;
        RECT 2475.785 145.695 2476.115 145.710 ;
        RECT 2567.785 145.695 2568.115 145.710 ;
        RECT 2668.985 145.695 2669.315 145.710 ;
        RECT 2762.365 145.695 2762.695 145.710 ;
        RECT 1917.590 145.030 1918.810 145.330 ;
        RECT 2863.350 145.330 2863.650 146.390 ;
        RECT 2916.710 146.390 2924.800 146.690 ;
        RECT 2916.710 145.330 2917.010 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
        RECT 2863.350 145.030 2917.010 145.330 ;
        RECT 1448.605 145.015 1448.935 145.030 ;
      LAYER via3 ;
        RECT 1158.580 1996.660 1158.900 1996.980 ;
        RECT 1158.580 145.020 1158.900 145.340 ;
      LAYER met4 ;
        RECT 1158.575 1996.655 1158.905 1996.985 ;
        RECT 1158.590 145.345 1158.890 1996.655 ;
        RECT 1158.575 145.015 1158.905 145.345 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1240.690 2491.080 1241.010 2491.140 ;
        RECT 2900.830 2491.080 2901.150 2491.140 ;
        RECT 1240.690 2490.940 2901.150 2491.080 ;
        RECT 1240.690 2490.880 1241.010 2490.940 ;
        RECT 2900.830 2490.880 2901.150 2490.940 ;
        RECT 1235.170 2009.640 1235.490 2009.700 ;
        RECT 1240.690 2009.640 1241.010 2009.700 ;
        RECT 1235.170 2009.500 1241.010 2009.640 ;
        RECT 1235.170 2009.440 1235.490 2009.500 ;
        RECT 1240.690 2009.440 1241.010 2009.500 ;
      LAYER via ;
        RECT 1240.720 2490.880 1240.980 2491.140 ;
        RECT 2900.860 2490.880 2901.120 2491.140 ;
        RECT 1235.200 2009.440 1235.460 2009.700 ;
        RECT 1240.720 2009.440 1240.980 2009.700 ;
      LAYER met2 ;
        RECT 2900.850 2493.035 2901.130 2493.405 ;
        RECT 2900.920 2491.170 2901.060 2493.035 ;
        RECT 1240.720 2490.850 1240.980 2491.170 ;
        RECT 2900.860 2490.850 2901.120 2491.170 ;
        RECT 1240.780 2009.730 1240.920 2490.850 ;
        RECT 1235.200 2009.410 1235.460 2009.730 ;
        RECT 1240.720 2009.410 1240.980 2009.730 ;
        RECT 1235.260 2000.000 1235.400 2009.410 ;
        RECT 1235.100 1999.540 1235.400 2000.000 ;
        RECT 1235.100 1996.000 1235.380 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2493.080 2901.130 2493.360 ;
      LAYER met3 ;
        RECT 2900.825 2493.370 2901.155 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.825 2493.070 2924.800 2493.370 ;
        RECT 2900.825 2493.055 2901.155 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1247.590 2725.680 1247.910 2725.740 ;
        RECT 2900.830 2725.680 2901.150 2725.740 ;
        RECT 1247.590 2725.540 2901.150 2725.680 ;
        RECT 1247.590 2725.480 1247.910 2725.540 ;
        RECT 2900.830 2725.480 2901.150 2725.540 ;
        RECT 1242.990 2010.660 1243.310 2010.720 ;
        RECT 1247.590 2010.660 1247.910 2010.720 ;
        RECT 1242.990 2010.520 1247.910 2010.660 ;
        RECT 1242.990 2010.460 1243.310 2010.520 ;
        RECT 1247.590 2010.460 1247.910 2010.520 ;
      LAYER via ;
        RECT 1247.620 2725.480 1247.880 2725.740 ;
        RECT 2900.860 2725.480 2901.120 2725.740 ;
        RECT 1243.020 2010.460 1243.280 2010.720 ;
        RECT 1247.620 2010.460 1247.880 2010.720 ;
      LAYER met2 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2725.770 2901.060 2727.635 ;
        RECT 1247.620 2725.450 1247.880 2725.770 ;
        RECT 2900.860 2725.450 2901.120 2725.770 ;
        RECT 1247.680 2010.750 1247.820 2725.450 ;
        RECT 1243.020 2010.430 1243.280 2010.750 ;
        RECT 1247.620 2010.430 1247.880 2010.750 ;
        RECT 1243.080 2000.000 1243.220 2010.430 ;
        RECT 1242.920 1999.540 1243.220 2000.000 ;
        RECT 1242.920 1996.000 1243.200 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
      LAYER met3 ;
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1254.950 2960.280 1255.270 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 1254.950 2960.140 2901.150 2960.280 ;
        RECT 1254.950 2960.080 1255.270 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
        RECT 1250.810 2010.660 1251.130 2010.720 ;
        RECT 1254.950 2010.660 1255.270 2010.720 ;
        RECT 1250.810 2010.520 1255.270 2010.660 ;
        RECT 1250.810 2010.460 1251.130 2010.520 ;
        RECT 1254.950 2010.460 1255.270 2010.520 ;
      LAYER via ;
        RECT 1254.980 2960.080 1255.240 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
        RECT 1250.840 2010.460 1251.100 2010.720 ;
        RECT 1254.980 2010.460 1255.240 2010.720 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 1254.980 2960.050 1255.240 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 1255.040 2010.750 1255.180 2960.050 ;
        RECT 1250.840 2010.430 1251.100 2010.750 ;
        RECT 1254.980 2010.430 1255.240 2010.750 ;
        RECT 1250.900 2000.000 1251.040 2010.430 ;
        RECT 1250.740 1999.540 1251.040 2000.000 ;
        RECT 1250.740 1996.000 1251.020 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
      LAYER met3 ;
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1261.390 3194.880 1261.710 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 1261.390 3194.740 2901.150 3194.880 ;
        RECT 1261.390 3194.680 1261.710 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
      LAYER via ;
        RECT 1261.420 3194.680 1261.680 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 1261.420 3194.650 1261.680 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 1261.480 2001.650 1261.620 3194.650 ;
        RECT 1261.020 2001.510 1261.620 2001.650 ;
        RECT 1258.560 1998.930 1258.840 2000.000 ;
        RECT 1261.020 1998.930 1261.160 2001.510 ;
        RECT 1258.560 1998.790 1261.160 1998.930 ;
        RECT 1258.560 1996.000 1258.840 1998.790 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1497.460 3429.680 1506.340 3429.820 ;
        RECT 1268.290 3429.480 1268.610 3429.540 ;
        RECT 1497.460 3429.480 1497.600 3429.680 ;
        RECT 1268.290 3429.340 1497.600 3429.480 ;
        RECT 1506.200 3429.480 1506.340 3429.680 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 1506.200 3429.340 2901.150 3429.480 ;
        RECT 1268.290 3429.280 1268.610 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 1268.320 3429.280 1268.580 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 1268.320 3429.250 1268.580 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 1266.380 1999.610 1266.660 2000.000 ;
        RECT 1268.380 1999.610 1268.520 3429.250 ;
        RECT 1266.380 1999.470 1268.520 1999.610 ;
        RECT 1266.380 1996.000 1266.660 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1275.650 3501.900 1275.970 3501.960 ;
        RECT 2717.290 3501.900 2717.610 3501.960 ;
        RECT 1275.650 3501.760 2717.610 3501.900 ;
        RECT 1275.650 3501.700 1275.970 3501.760 ;
        RECT 2717.290 3501.700 2717.610 3501.760 ;
      LAYER via ;
        RECT 1275.680 3501.700 1275.940 3501.960 ;
        RECT 2717.320 3501.700 2717.580 3501.960 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.990 2717.520 3517.600 ;
        RECT 1275.680 3501.670 1275.940 3501.990 ;
        RECT 2717.320 3501.670 2717.580 3501.990 ;
        RECT 1274.200 1999.610 1274.480 2000.000 ;
        RECT 1275.740 1999.610 1275.880 3501.670 ;
        RECT 1274.200 1999.470 1275.880 1999.610 ;
        RECT 1274.200 1996.000 1274.480 1999.470 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1282.550 3503.260 1282.870 3503.320 ;
        RECT 2392.530 3503.260 2392.850 3503.320 ;
        RECT 1282.550 3503.120 2392.850 3503.260 ;
        RECT 1282.550 3503.060 1282.870 3503.120 ;
        RECT 2392.530 3503.060 2392.850 3503.120 ;
      LAYER via ;
        RECT 1282.580 3503.060 1282.840 3503.320 ;
        RECT 2392.560 3503.060 2392.820 3503.320 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3503.350 2392.760 3517.600 ;
        RECT 1282.580 3503.030 1282.840 3503.350 ;
        RECT 2392.560 3503.030 2392.820 3503.350 ;
        RECT 1282.020 1999.610 1282.300 2000.000 ;
        RECT 1282.640 1999.610 1282.780 3503.030 ;
        RECT 1282.020 1999.470 1282.780 1999.610 ;
        RECT 1282.020 1996.000 1282.300 1999.470 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1296.350 3504.620 1296.670 3504.680 ;
        RECT 2068.230 3504.620 2068.550 3504.680 ;
        RECT 1296.350 3504.480 2068.550 3504.620 ;
        RECT 1296.350 3504.420 1296.670 3504.480 ;
        RECT 2068.230 3504.420 2068.550 3504.480 ;
        RECT 1292.210 2038.880 1292.530 2038.940 ;
        RECT 1296.350 2038.880 1296.670 2038.940 ;
        RECT 1292.210 2038.740 1296.670 2038.880 ;
        RECT 1292.210 2038.680 1292.530 2038.740 ;
        RECT 1296.350 2038.680 1296.670 2038.740 ;
      LAYER via ;
        RECT 1296.380 3504.420 1296.640 3504.680 ;
        RECT 2068.260 3504.420 2068.520 3504.680 ;
        RECT 1292.240 2038.680 1292.500 2038.940 ;
        RECT 1296.380 2038.680 1296.640 2038.940 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3504.710 2068.460 3517.600 ;
        RECT 1296.380 3504.390 1296.640 3504.710 ;
        RECT 2068.260 3504.390 2068.520 3504.710 ;
        RECT 1296.440 2038.970 1296.580 3504.390 ;
        RECT 1292.240 2038.650 1292.500 2038.970 ;
        RECT 1296.380 2038.650 1296.640 2038.970 ;
        RECT 1290.300 1999.610 1290.580 2000.000 ;
        RECT 1292.300 1999.610 1292.440 2038.650 ;
        RECT 1290.300 1999.470 1292.440 1999.610 ;
        RECT 1290.300 1996.000 1290.580 1999.470 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1303.250 3500.540 1303.570 3500.600 ;
        RECT 1743.930 3500.540 1744.250 3500.600 ;
        RECT 1303.250 3500.400 1744.250 3500.540 ;
        RECT 1303.250 3500.340 1303.570 3500.400 ;
        RECT 1743.930 3500.340 1744.250 3500.400 ;
        RECT 1298.190 2010.320 1298.510 2010.380 ;
        RECT 1303.250 2010.320 1303.570 2010.380 ;
        RECT 1298.190 2010.180 1303.570 2010.320 ;
        RECT 1298.190 2010.120 1298.510 2010.180 ;
        RECT 1303.250 2010.120 1303.570 2010.180 ;
      LAYER via ;
        RECT 1303.280 3500.340 1303.540 3500.600 ;
        RECT 1743.960 3500.340 1744.220 3500.600 ;
        RECT 1298.220 2010.120 1298.480 2010.380 ;
        RECT 1303.280 2010.120 1303.540 2010.380 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3500.630 1744.160 3517.600 ;
        RECT 1303.280 3500.310 1303.540 3500.630 ;
        RECT 1743.960 3500.310 1744.220 3500.630 ;
        RECT 1303.340 2010.410 1303.480 3500.310 ;
        RECT 1298.220 2010.090 1298.480 2010.410 ;
        RECT 1303.280 2010.090 1303.540 2010.410 ;
        RECT 1298.280 2000.000 1298.420 2010.090 ;
        RECT 1298.120 1999.540 1298.420 2000.000 ;
        RECT 1298.120 1996.000 1298.400 1999.540 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1310.610 3499.520 1310.930 3499.580 ;
        RECT 1419.170 3499.520 1419.490 3499.580 ;
        RECT 1310.610 3499.380 1419.490 3499.520 ;
        RECT 1310.610 3499.320 1310.930 3499.380 ;
        RECT 1419.170 3499.320 1419.490 3499.380 ;
        RECT 1306.010 2010.320 1306.330 2010.380 ;
        RECT 1310.610 2010.320 1310.930 2010.380 ;
        RECT 1306.010 2010.180 1310.930 2010.320 ;
        RECT 1306.010 2010.120 1306.330 2010.180 ;
        RECT 1310.610 2010.120 1310.930 2010.180 ;
      LAYER via ;
        RECT 1310.640 3499.320 1310.900 3499.580 ;
        RECT 1419.200 3499.320 1419.460 3499.580 ;
        RECT 1306.040 2010.120 1306.300 2010.380 ;
        RECT 1310.640 2010.120 1310.900 2010.380 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3499.610 1419.400 3517.600 ;
        RECT 1310.640 3499.290 1310.900 3499.610 ;
        RECT 1419.200 3499.290 1419.460 3499.610 ;
        RECT 1310.700 2010.410 1310.840 3499.290 ;
        RECT 1306.040 2010.090 1306.300 2010.410 ;
        RECT 1310.640 2010.090 1310.900 2010.410 ;
        RECT 1306.100 2000.000 1306.240 2010.090 ;
        RECT 1305.940 1999.540 1306.240 2000.000 ;
        RECT 1305.940 1996.000 1306.220 1999.540 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2766.510 380.700 2766.830 380.760 ;
        RECT 2772.950 380.700 2773.270 380.760 ;
        RECT 2766.510 380.560 2773.270 380.700 ;
        RECT 2766.510 380.500 2766.830 380.560 ;
        RECT 2772.950 380.500 2773.270 380.560 ;
        RECT 2186.910 380.360 2187.230 380.420 ;
        RECT 2221.410 380.360 2221.730 380.420 ;
        RECT 2186.910 380.220 2221.730 380.360 ;
        RECT 2186.910 380.160 2187.230 380.220 ;
        RECT 2221.410 380.160 2221.730 380.220 ;
        RECT 2511.210 380.360 2511.530 380.420 ;
        RECT 2552.610 380.360 2552.930 380.420 ;
        RECT 2511.210 380.220 2552.930 380.360 ;
        RECT 2511.210 380.160 2511.530 380.220 ;
        RECT 2552.610 380.160 2552.930 380.220 ;
        RECT 2669.910 380.360 2670.230 380.420 ;
        RECT 2704.410 380.360 2704.730 380.420 ;
        RECT 2669.910 380.220 2704.730 380.360 ;
        RECT 2669.910 380.160 2670.230 380.220 ;
        RECT 2704.410 380.160 2704.730 380.220 ;
        RECT 1545.670 380.020 1545.990 380.080 ;
        RECT 1569.590 380.020 1569.910 380.080 ;
        RECT 1545.670 379.880 1569.910 380.020 ;
        RECT 1545.670 379.820 1545.990 379.880 ;
        RECT 1569.590 379.820 1569.910 379.880 ;
      LAYER via ;
        RECT 2766.540 380.500 2766.800 380.760 ;
        RECT 2772.980 380.500 2773.240 380.760 ;
        RECT 2186.940 380.160 2187.200 380.420 ;
        RECT 2221.440 380.160 2221.700 380.420 ;
        RECT 2511.240 380.160 2511.500 380.420 ;
        RECT 2552.640 380.160 2552.900 380.420 ;
        RECT 2669.940 380.160 2670.200 380.420 ;
        RECT 2704.440 380.160 2704.700 380.420 ;
        RECT 1545.700 379.820 1545.960 380.080 ;
        RECT 1569.620 379.820 1569.880 380.080 ;
      LAYER met2 ;
        RECT 1163.800 1996.890 1164.080 2000.000 ;
        RECT 1164.810 1996.890 1165.090 1997.005 ;
        RECT 1163.800 1996.750 1165.090 1996.890 ;
        RECT 1163.800 1996.000 1164.080 1996.750 ;
        RECT 1164.810 1996.635 1165.090 1996.750 ;
        RECT 2607.830 382.315 2608.110 382.685 ;
        RECT 1642.290 381.210 1642.570 381.325 ;
        RECT 1642.290 381.070 1642.960 381.210 ;
        RECT 1642.290 380.955 1642.570 381.070 ;
        RECT 1510.730 380.275 1511.010 380.645 ;
        RECT 1569.610 380.275 1569.890 380.645 ;
        RECT 1617.910 380.275 1618.190 380.645 ;
        RECT 1510.800 378.605 1510.940 380.275 ;
        RECT 1569.680 380.110 1569.820 380.275 ;
        RECT 1545.700 379.965 1545.960 380.110 ;
        RECT 1545.690 379.595 1545.970 379.965 ;
        RECT 1569.620 379.790 1569.880 380.110 ;
        RECT 1617.980 379.285 1618.120 380.275 ;
        RECT 1642.820 379.285 1642.960 381.070 ;
        RECT 2552.630 380.955 2552.910 381.325 ;
        RECT 2076.530 380.275 2076.810 380.645 ;
        RECT 2186.930 380.275 2187.210 380.645 ;
        RECT 2283.530 380.530 2283.810 380.645 ;
        RECT 2284.450 380.530 2284.730 380.645 ;
        RECT 2076.600 379.965 2076.740 380.275 ;
        RECT 2186.940 380.130 2187.200 380.275 ;
        RECT 2221.440 380.130 2221.700 380.450 ;
        RECT 2283.530 380.390 2284.730 380.530 ;
        RECT 2283.530 380.275 2283.810 380.390 ;
        RECT 2284.450 380.275 2284.730 380.390 ;
        RECT 2414.630 380.275 2414.910 380.645 ;
        RECT 2552.700 380.450 2552.840 380.955 ;
        RECT 2221.500 379.965 2221.640 380.130 ;
        RECT 2414.700 379.965 2414.840 380.275 ;
        RECT 2511.240 380.130 2511.500 380.450 ;
        RECT 2552.640 380.130 2552.900 380.450 ;
        RECT 2076.530 379.595 2076.810 379.965 ;
        RECT 2221.430 379.595 2221.710 379.965 ;
        RECT 2414.630 379.595 2414.910 379.965 ;
        RECT 2511.300 379.285 2511.440 380.130 ;
        RECT 2607.900 379.965 2608.040 382.315 ;
        RECT 2766.540 380.645 2766.800 380.790 ;
        RECT 2772.980 380.645 2773.240 380.790 ;
        RECT 2669.930 380.275 2670.210 380.645 ;
        RECT 2669.940 380.130 2670.200 380.275 ;
        RECT 2704.440 380.130 2704.700 380.450 ;
        RECT 2766.530 380.275 2766.810 380.645 ;
        RECT 2772.970 380.275 2773.250 380.645 ;
        RECT 2704.500 379.965 2704.640 380.130 ;
        RECT 2607.830 379.595 2608.110 379.965 ;
        RECT 2704.430 379.595 2704.710 379.965 ;
        RECT 1617.910 378.915 1618.190 379.285 ;
        RECT 1642.750 378.915 1643.030 379.285 ;
        RECT 2511.230 378.915 2511.510 379.285 ;
        RECT 1510.730 378.235 1511.010 378.605 ;
      LAYER via2 ;
        RECT 1164.810 1996.680 1165.090 1996.960 ;
        RECT 2607.830 382.360 2608.110 382.640 ;
        RECT 1642.290 381.000 1642.570 381.280 ;
        RECT 1510.730 380.320 1511.010 380.600 ;
        RECT 1569.610 380.320 1569.890 380.600 ;
        RECT 1617.910 380.320 1618.190 380.600 ;
        RECT 1545.690 379.640 1545.970 379.920 ;
        RECT 2552.630 381.000 2552.910 381.280 ;
        RECT 2076.530 380.320 2076.810 380.600 ;
        RECT 2186.930 380.320 2187.210 380.600 ;
        RECT 2283.530 380.320 2283.810 380.600 ;
        RECT 2284.450 380.320 2284.730 380.600 ;
        RECT 2414.630 380.320 2414.910 380.600 ;
        RECT 2076.530 379.640 2076.810 379.920 ;
        RECT 2221.430 379.640 2221.710 379.920 ;
        RECT 2414.630 379.640 2414.910 379.920 ;
        RECT 2669.930 380.320 2670.210 380.600 ;
        RECT 2766.530 380.320 2766.810 380.600 ;
        RECT 2772.970 380.320 2773.250 380.600 ;
        RECT 2607.830 379.640 2608.110 379.920 ;
        RECT 2704.430 379.640 2704.710 379.920 ;
        RECT 1617.910 378.960 1618.190 379.240 ;
        RECT 1642.750 378.960 1643.030 379.240 ;
        RECT 2511.230 378.960 2511.510 379.240 ;
        RECT 1510.730 378.280 1511.010 378.560 ;
      LAYER met3 ;
        RECT 1164.785 1996.980 1165.115 1996.985 ;
        RECT 1164.785 1996.970 1165.370 1996.980 ;
        RECT 1164.785 1996.670 1165.570 1996.970 ;
        RECT 1164.785 1996.660 1165.370 1996.670 ;
        RECT 1164.785 1996.655 1165.115 1996.660 ;
        RECT 2607.805 382.650 2608.135 382.665 ;
        RECT 2559.750 382.350 2608.135 382.650 ;
        RECT 1164.990 381.290 1165.370 381.300 ;
        RECT 1642.265 381.290 1642.595 381.305 ;
        RECT 1164.990 380.990 1172.690 381.290 ;
        RECT 1164.990 380.980 1165.370 380.990 ;
        RECT 1172.390 379.930 1172.690 380.990 ;
        RECT 1173.310 380.990 1231.570 381.290 ;
        RECT 1173.310 379.930 1173.610 380.990 ;
        RECT 1172.390 379.630 1173.610 379.930 ;
        RECT 1231.270 379.930 1231.570 380.990 ;
        RECT 1641.590 380.990 1642.595 381.290 ;
        RECT 1510.705 380.610 1511.035 380.625 ;
        RECT 1463.110 380.310 1511.035 380.610 ;
        RECT 1463.110 379.930 1463.410 380.310 ;
        RECT 1510.705 380.295 1511.035 380.310 ;
        RECT 1569.585 380.610 1569.915 380.625 ;
        RECT 1593.710 380.610 1594.090 380.620 ;
        RECT 1569.585 380.310 1594.090 380.610 ;
        RECT 1569.585 380.295 1569.915 380.310 ;
        RECT 1593.710 380.300 1594.090 380.310 ;
        RECT 1617.885 380.610 1618.215 380.625 ;
        RECT 1641.590 380.610 1641.890 380.990 ;
        RECT 1642.265 380.975 1642.595 380.990 ;
        RECT 1690.310 381.290 1690.690 381.300 ;
        RECT 2552.605 381.290 2552.935 381.305 ;
        RECT 2559.750 381.290 2560.050 382.350 ;
        RECT 2607.805 382.335 2608.135 382.350 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 1690.310 380.990 1773.450 381.290 ;
        RECT 1690.310 380.980 1690.690 380.990 ;
        RECT 1617.885 380.310 1641.890 380.610 ;
        RECT 1773.150 380.610 1773.450 380.990 ;
        RECT 1821.910 380.990 1870.050 381.290 ;
        RECT 1773.150 380.310 1821.290 380.610 ;
        RECT 1617.885 380.295 1618.215 380.310 ;
        RECT 1545.665 379.930 1545.995 379.945 ;
        RECT 1690.310 379.930 1690.690 379.940 ;
        RECT 1231.270 379.630 1463.410 379.930 ;
        RECT 1544.990 379.630 1545.995 379.930 ;
        RECT 1510.705 378.570 1511.035 378.585 ;
        RECT 1544.990 378.570 1545.290 379.630 ;
        RECT 1545.665 379.615 1545.995 379.630 ;
        RECT 1657.230 379.630 1690.690 379.930 ;
        RECT 1820.990 379.930 1821.290 380.310 ;
        RECT 1821.910 379.930 1822.210 380.990 ;
        RECT 1869.750 380.610 1870.050 380.990 ;
        RECT 1918.510 380.990 2029.210 381.290 ;
        RECT 1869.750 380.310 1917.890 380.610 ;
        RECT 1820.990 379.630 1822.210 379.930 ;
        RECT 1917.590 379.930 1917.890 380.310 ;
        RECT 1918.510 379.930 1918.810 380.990 ;
        RECT 2028.910 380.610 2029.210 380.990 ;
        RECT 2552.605 380.990 2560.050 381.290 ;
        RECT 2916.710 380.990 2924.800 381.290 ;
        RECT 2552.605 380.975 2552.935 380.990 ;
        RECT 2076.505 380.610 2076.835 380.625 ;
        RECT 2186.905 380.610 2187.235 380.625 ;
        RECT 2283.505 380.610 2283.835 380.625 ;
        RECT 2028.910 380.310 2076.835 380.610 ;
        RECT 2076.505 380.295 2076.835 380.310 ;
        RECT 2139.310 380.310 2187.235 380.610 ;
        RECT 1917.590 379.630 1918.810 379.930 ;
        RECT 2076.505 379.930 2076.835 379.945 ;
        RECT 2139.310 379.930 2139.610 380.310 ;
        RECT 2186.905 380.295 2187.235 380.310 ;
        RECT 2235.910 380.310 2283.835 380.610 ;
        RECT 2076.505 379.630 2139.610 379.930 ;
        RECT 2221.405 379.930 2221.735 379.945 ;
        RECT 2235.910 379.930 2236.210 380.310 ;
        RECT 2283.505 380.295 2283.835 380.310 ;
        RECT 2284.425 380.610 2284.755 380.625 ;
        RECT 2414.605 380.610 2414.935 380.625 ;
        RECT 2463.110 380.610 2463.490 380.620 ;
        RECT 2669.905 380.610 2670.235 380.625 ;
        RECT 2766.505 380.610 2766.835 380.625 ;
        RECT 2284.425 380.310 2331.890 380.610 ;
        RECT 2284.425 380.295 2284.755 380.310 ;
        RECT 2221.405 379.630 2236.210 379.930 ;
        RECT 2331.590 379.930 2331.890 380.310 ;
        RECT 2332.510 380.310 2414.935 380.610 ;
        RECT 2332.510 379.930 2332.810 380.310 ;
        RECT 2414.605 380.295 2414.935 380.310 ;
        RECT 2415.310 380.310 2463.490 380.610 ;
        RECT 2331.590 379.630 2332.810 379.930 ;
        RECT 2414.605 379.930 2414.935 379.945 ;
        RECT 2415.310 379.930 2415.610 380.310 ;
        RECT 2463.110 380.300 2463.490 380.310 ;
        RECT 2622.310 380.310 2670.235 380.610 ;
        RECT 2414.605 379.630 2415.610 379.930 ;
        RECT 2607.805 379.930 2608.135 379.945 ;
        RECT 2622.310 379.930 2622.610 380.310 ;
        RECT 2669.905 380.295 2670.235 380.310 ;
        RECT 2718.910 380.310 2766.835 380.610 ;
        RECT 2607.805 379.630 2622.610 379.930 ;
        RECT 2704.405 379.930 2704.735 379.945 ;
        RECT 2718.910 379.930 2719.210 380.310 ;
        RECT 2766.505 380.295 2766.835 380.310 ;
        RECT 2772.945 380.610 2773.275 380.625 ;
        RECT 2916.710 380.610 2917.010 380.990 ;
        RECT 2772.945 380.310 2814.890 380.610 ;
        RECT 2772.945 380.295 2773.275 380.310 ;
        RECT 2704.405 379.630 2719.210 379.930 ;
        RECT 2814.590 379.930 2814.890 380.310 ;
        RECT 2884.510 380.310 2917.010 380.610 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
        RECT 2884.510 379.930 2884.810 380.310 ;
        RECT 2814.590 379.630 2884.810 379.930 ;
        RECT 1593.710 379.250 1594.090 379.260 ;
        RECT 1617.885 379.250 1618.215 379.265 ;
        RECT 1593.710 378.950 1618.215 379.250 ;
        RECT 1593.710 378.940 1594.090 378.950 ;
        RECT 1617.885 378.935 1618.215 378.950 ;
        RECT 1642.725 379.250 1643.055 379.265 ;
        RECT 1657.230 379.250 1657.530 379.630 ;
        RECT 1690.310 379.620 1690.690 379.630 ;
        RECT 2076.505 379.615 2076.835 379.630 ;
        RECT 2221.405 379.615 2221.735 379.630 ;
        RECT 2414.605 379.615 2414.935 379.630 ;
        RECT 2607.805 379.615 2608.135 379.630 ;
        RECT 2704.405 379.615 2704.735 379.630 ;
        RECT 1642.725 378.950 1657.530 379.250 ;
        RECT 2463.110 379.250 2463.490 379.260 ;
        RECT 2511.205 379.250 2511.535 379.265 ;
        RECT 2463.110 378.950 2511.535 379.250 ;
        RECT 1642.725 378.935 1643.055 378.950 ;
        RECT 2463.110 378.940 2463.490 378.950 ;
        RECT 2511.205 378.935 2511.535 378.950 ;
        RECT 1510.705 378.270 1545.290 378.570 ;
        RECT 1510.705 378.255 1511.035 378.270 ;
      LAYER via3 ;
        RECT 1165.020 1996.660 1165.340 1996.980 ;
        RECT 1165.020 380.980 1165.340 381.300 ;
        RECT 1593.740 380.300 1594.060 380.620 ;
        RECT 1690.340 380.980 1690.660 381.300 ;
        RECT 1593.740 378.940 1594.060 379.260 ;
        RECT 1690.340 379.620 1690.660 379.940 ;
        RECT 2463.140 380.300 2463.460 380.620 ;
        RECT 2463.140 378.940 2463.460 379.260 ;
      LAYER met4 ;
        RECT 1165.015 1996.655 1165.345 1996.985 ;
        RECT 1165.030 381.305 1165.330 1996.655 ;
        RECT 1165.015 380.975 1165.345 381.305 ;
        RECT 1690.335 380.975 1690.665 381.305 ;
        RECT 1593.735 380.295 1594.065 380.625 ;
        RECT 1593.750 379.265 1594.050 380.295 ;
        RECT 1690.350 379.945 1690.650 380.975 ;
        RECT 2463.135 380.295 2463.465 380.625 ;
        RECT 1690.335 379.615 1690.665 379.945 ;
        RECT 2463.150 379.265 2463.450 380.295 ;
        RECT 1593.735 378.935 1594.065 379.265 ;
        RECT 2463.135 378.935 2463.465 379.265 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1095.405 3429.325 1095.575 3477.435 ;
        RECT 1094.945 3332.765 1095.115 3380.875 ;
        RECT 1096.325 3236.205 1096.495 3284.315 ;
        RECT 1096.785 3084.225 1096.955 3132.675 ;
        RECT 1095.405 3043.425 1095.575 3057.195 ;
        RECT 1096.325 3007.725 1096.495 3042.915 ;
        RECT 1095.865 2946.525 1096.035 2994.635 ;
        RECT 1094.485 2849.625 1094.655 2898.075 ;
        RECT 1094.485 2753.065 1094.655 2767.175 ;
        RECT 1095.405 2525.265 1095.575 2552.975 ;
        RECT 1094.945 2221.985 1095.115 2270.095 ;
      LAYER mcon ;
        RECT 1095.405 3477.265 1095.575 3477.435 ;
        RECT 1094.945 3380.705 1095.115 3380.875 ;
        RECT 1096.325 3284.145 1096.495 3284.315 ;
        RECT 1096.785 3132.505 1096.955 3132.675 ;
        RECT 1095.405 3057.025 1095.575 3057.195 ;
        RECT 1096.325 3042.745 1096.495 3042.915 ;
        RECT 1095.865 2994.465 1096.035 2994.635 ;
        RECT 1094.485 2897.905 1094.655 2898.075 ;
        RECT 1094.485 2767.005 1094.655 2767.175 ;
        RECT 1095.405 2552.805 1095.575 2552.975 ;
        RECT 1094.945 2269.925 1095.115 2270.095 ;
      LAYER met1 ;
        RECT 1095.345 3477.420 1095.635 3477.465 ;
        RECT 1095.790 3477.420 1096.110 3477.480 ;
        RECT 1095.345 3477.280 1096.110 3477.420 ;
        RECT 1095.345 3477.235 1095.635 3477.280 ;
        RECT 1095.790 3477.220 1096.110 3477.280 ;
        RECT 1095.330 3429.480 1095.650 3429.540 ;
        RECT 1095.135 3429.340 1095.650 3429.480 ;
        RECT 1095.330 3429.280 1095.650 3429.340 ;
        RECT 1094.870 3380.860 1095.190 3380.920 ;
        RECT 1094.675 3380.720 1095.190 3380.860 ;
        RECT 1094.870 3380.660 1095.190 3380.720 ;
        RECT 1094.885 3332.920 1095.175 3332.965 ;
        RECT 1095.330 3332.920 1095.650 3332.980 ;
        RECT 1094.885 3332.780 1095.650 3332.920 ;
        RECT 1094.885 3332.735 1095.175 3332.780 ;
        RECT 1095.330 3332.720 1095.650 3332.780 ;
        RECT 1095.790 3298.240 1096.110 3298.300 ;
        RECT 1096.710 3298.240 1097.030 3298.300 ;
        RECT 1095.790 3298.100 1097.030 3298.240 ;
        RECT 1095.790 3298.040 1096.110 3298.100 ;
        RECT 1096.710 3298.040 1097.030 3298.100 ;
        RECT 1096.265 3284.300 1096.555 3284.345 ;
        RECT 1096.710 3284.300 1097.030 3284.360 ;
        RECT 1096.265 3284.160 1097.030 3284.300 ;
        RECT 1096.265 3284.115 1096.555 3284.160 ;
        RECT 1096.710 3284.100 1097.030 3284.160 ;
        RECT 1096.250 3236.360 1096.570 3236.420 ;
        RECT 1096.055 3236.220 1096.570 3236.360 ;
        RECT 1096.250 3236.160 1096.570 3236.220 ;
        RECT 1096.250 3202.020 1096.570 3202.080 ;
        RECT 1095.420 3201.880 1096.570 3202.020 ;
        RECT 1095.420 3201.400 1095.560 3201.880 ;
        RECT 1096.250 3201.820 1096.570 3201.880 ;
        RECT 1095.330 3201.140 1095.650 3201.400 ;
        RECT 1095.330 3187.740 1095.650 3187.800 ;
        RECT 1095.790 3187.740 1096.110 3187.800 ;
        RECT 1095.330 3187.600 1096.110 3187.740 ;
        RECT 1095.330 3187.540 1095.650 3187.600 ;
        RECT 1095.790 3187.540 1096.110 3187.600 ;
        RECT 1096.710 3132.660 1097.030 3132.720 ;
        RECT 1096.515 3132.520 1097.030 3132.660 ;
        RECT 1096.710 3132.460 1097.030 3132.520 ;
        RECT 1096.710 3084.380 1097.030 3084.440 ;
        RECT 1096.515 3084.240 1097.030 3084.380 ;
        RECT 1096.710 3084.180 1097.030 3084.240 ;
        RECT 1095.345 3057.180 1095.635 3057.225 ;
        RECT 1096.710 3057.180 1097.030 3057.240 ;
        RECT 1095.345 3057.040 1097.030 3057.180 ;
        RECT 1095.345 3056.995 1095.635 3057.040 ;
        RECT 1096.710 3056.980 1097.030 3057.040 ;
        RECT 1095.330 3043.580 1095.650 3043.640 ;
        RECT 1095.135 3043.440 1095.650 3043.580 ;
        RECT 1095.330 3043.380 1095.650 3043.440 ;
        RECT 1095.330 3042.900 1095.650 3042.960 ;
        RECT 1096.265 3042.900 1096.555 3042.945 ;
        RECT 1095.330 3042.760 1096.555 3042.900 ;
        RECT 1095.330 3042.700 1095.650 3042.760 ;
        RECT 1096.265 3042.715 1096.555 3042.760 ;
        RECT 1096.250 3007.880 1096.570 3007.940 ;
        RECT 1096.055 3007.740 1096.570 3007.880 ;
        RECT 1096.250 3007.680 1096.570 3007.740 ;
        RECT 1095.805 2994.620 1096.095 2994.665 ;
        RECT 1096.250 2994.620 1096.570 2994.680 ;
        RECT 1095.805 2994.480 1096.570 2994.620 ;
        RECT 1095.805 2994.435 1096.095 2994.480 ;
        RECT 1096.250 2994.420 1096.570 2994.480 ;
        RECT 1095.790 2946.680 1096.110 2946.740 ;
        RECT 1095.595 2946.540 1096.110 2946.680 ;
        RECT 1095.790 2946.480 1096.110 2946.540 ;
        RECT 1094.870 2912.000 1095.190 2912.060 ;
        RECT 1095.790 2912.000 1096.110 2912.060 ;
        RECT 1094.870 2911.860 1096.110 2912.000 ;
        RECT 1094.870 2911.800 1095.190 2911.860 ;
        RECT 1095.790 2911.800 1096.110 2911.860 ;
        RECT 1094.425 2898.060 1094.715 2898.105 ;
        RECT 1094.870 2898.060 1095.190 2898.120 ;
        RECT 1094.425 2897.920 1095.190 2898.060 ;
        RECT 1094.425 2897.875 1094.715 2897.920 ;
        RECT 1094.870 2897.860 1095.190 2897.920 ;
        RECT 1094.410 2849.780 1094.730 2849.840 ;
        RECT 1094.215 2849.640 1094.730 2849.780 ;
        RECT 1094.410 2849.580 1094.730 2849.640 ;
        RECT 1094.410 2815.240 1094.730 2815.500 ;
        RECT 1094.500 2814.760 1094.640 2815.240 ;
        RECT 1094.870 2814.760 1095.190 2814.820 ;
        RECT 1094.500 2814.620 1095.190 2814.760 ;
        RECT 1094.870 2814.560 1095.190 2814.620 ;
        RECT 1094.410 2767.160 1094.730 2767.220 ;
        RECT 1094.215 2767.020 1094.730 2767.160 ;
        RECT 1094.410 2766.960 1094.730 2767.020 ;
        RECT 1094.410 2753.220 1094.730 2753.280 ;
        RECT 1094.215 2753.080 1094.730 2753.220 ;
        RECT 1094.410 2753.020 1094.730 2753.080 ;
        RECT 1094.410 2718.680 1094.730 2718.940 ;
        RECT 1094.500 2718.200 1094.640 2718.680 ;
        RECT 1094.870 2718.200 1095.190 2718.260 ;
        RECT 1094.500 2718.060 1095.190 2718.200 ;
        RECT 1094.870 2718.000 1095.190 2718.060 ;
        RECT 1094.870 2621.640 1095.190 2621.700 ;
        RECT 1095.790 2621.640 1096.110 2621.700 ;
        RECT 1094.870 2621.500 1096.110 2621.640 ;
        RECT 1094.870 2621.440 1095.190 2621.500 ;
        RECT 1095.790 2621.440 1096.110 2621.500 ;
        RECT 1093.950 2573.360 1094.270 2573.420 ;
        RECT 1095.330 2573.360 1095.650 2573.420 ;
        RECT 1093.950 2573.220 1095.650 2573.360 ;
        RECT 1093.950 2573.160 1094.270 2573.220 ;
        RECT 1095.330 2573.160 1095.650 2573.220 ;
        RECT 1095.330 2552.960 1095.650 2553.020 ;
        RECT 1095.135 2552.820 1095.650 2552.960 ;
        RECT 1095.330 2552.760 1095.650 2552.820 ;
        RECT 1095.330 2525.420 1095.650 2525.480 ;
        RECT 1095.135 2525.280 1095.650 2525.420 ;
        RECT 1095.330 2525.220 1095.650 2525.280 ;
        RECT 1095.330 2463.540 1095.650 2463.600 ;
        RECT 1095.790 2463.540 1096.110 2463.600 ;
        RECT 1095.330 2463.400 1096.110 2463.540 ;
        RECT 1095.330 2463.340 1095.650 2463.400 ;
        RECT 1095.790 2463.340 1096.110 2463.400 ;
        RECT 1095.790 2429.000 1096.110 2429.260 ;
        RECT 1095.880 2428.520 1096.020 2429.000 ;
        RECT 1096.250 2428.520 1096.570 2428.580 ;
        RECT 1095.880 2428.380 1096.570 2428.520 ;
        RECT 1096.250 2428.320 1096.570 2428.380 ;
        RECT 1094.870 2332.100 1095.190 2332.360 ;
        RECT 1094.960 2331.620 1095.100 2332.100 ;
        RECT 1096.710 2331.620 1097.030 2331.680 ;
        RECT 1094.960 2331.480 1097.030 2331.620 ;
        RECT 1096.710 2331.420 1097.030 2331.480 ;
        RECT 1094.885 2270.080 1095.175 2270.125 ;
        RECT 1095.330 2270.080 1095.650 2270.140 ;
        RECT 1094.885 2269.940 1095.650 2270.080 ;
        RECT 1094.885 2269.895 1095.175 2269.940 ;
        RECT 1095.330 2269.880 1095.650 2269.940 ;
        RECT 1094.870 2222.140 1095.190 2222.200 ;
        RECT 1094.675 2222.000 1095.190 2222.140 ;
        RECT 1094.870 2221.940 1095.190 2222.000 ;
        RECT 1094.870 2173.520 1095.190 2173.580 ;
        RECT 1095.330 2173.520 1095.650 2173.580 ;
        RECT 1094.870 2173.380 1095.650 2173.520 ;
        RECT 1094.870 2173.320 1095.190 2173.380 ;
        RECT 1095.330 2173.320 1095.650 2173.380 ;
        RECT 1096.710 2011.000 1097.030 2011.060 ;
        RECT 1313.830 2011.000 1314.150 2011.060 ;
        RECT 1096.710 2010.860 1314.150 2011.000 ;
        RECT 1096.710 2010.800 1097.030 2010.860 ;
        RECT 1313.830 2010.800 1314.150 2010.860 ;
      LAYER via ;
        RECT 1095.820 3477.220 1096.080 3477.480 ;
        RECT 1095.360 3429.280 1095.620 3429.540 ;
        RECT 1094.900 3380.660 1095.160 3380.920 ;
        RECT 1095.360 3332.720 1095.620 3332.980 ;
        RECT 1095.820 3298.040 1096.080 3298.300 ;
        RECT 1096.740 3298.040 1097.000 3298.300 ;
        RECT 1096.740 3284.100 1097.000 3284.360 ;
        RECT 1096.280 3236.160 1096.540 3236.420 ;
        RECT 1096.280 3201.820 1096.540 3202.080 ;
        RECT 1095.360 3201.140 1095.620 3201.400 ;
        RECT 1095.360 3187.540 1095.620 3187.800 ;
        RECT 1095.820 3187.540 1096.080 3187.800 ;
        RECT 1096.740 3132.460 1097.000 3132.720 ;
        RECT 1096.740 3084.180 1097.000 3084.440 ;
        RECT 1096.740 3056.980 1097.000 3057.240 ;
        RECT 1095.360 3043.380 1095.620 3043.640 ;
        RECT 1095.360 3042.700 1095.620 3042.960 ;
        RECT 1096.280 3007.680 1096.540 3007.940 ;
        RECT 1096.280 2994.420 1096.540 2994.680 ;
        RECT 1095.820 2946.480 1096.080 2946.740 ;
        RECT 1094.900 2911.800 1095.160 2912.060 ;
        RECT 1095.820 2911.800 1096.080 2912.060 ;
        RECT 1094.900 2897.860 1095.160 2898.120 ;
        RECT 1094.440 2849.580 1094.700 2849.840 ;
        RECT 1094.440 2815.240 1094.700 2815.500 ;
        RECT 1094.900 2814.560 1095.160 2814.820 ;
        RECT 1094.440 2766.960 1094.700 2767.220 ;
        RECT 1094.440 2753.020 1094.700 2753.280 ;
        RECT 1094.440 2718.680 1094.700 2718.940 ;
        RECT 1094.900 2718.000 1095.160 2718.260 ;
        RECT 1094.900 2621.440 1095.160 2621.700 ;
        RECT 1095.820 2621.440 1096.080 2621.700 ;
        RECT 1093.980 2573.160 1094.240 2573.420 ;
        RECT 1095.360 2573.160 1095.620 2573.420 ;
        RECT 1095.360 2552.760 1095.620 2553.020 ;
        RECT 1095.360 2525.220 1095.620 2525.480 ;
        RECT 1095.360 2463.340 1095.620 2463.600 ;
        RECT 1095.820 2463.340 1096.080 2463.600 ;
        RECT 1095.820 2429.000 1096.080 2429.260 ;
        RECT 1096.280 2428.320 1096.540 2428.580 ;
        RECT 1094.900 2332.100 1095.160 2332.360 ;
        RECT 1096.740 2331.420 1097.000 2331.680 ;
        RECT 1095.360 2269.880 1095.620 2270.140 ;
        RECT 1094.900 2221.940 1095.160 2222.200 ;
        RECT 1094.900 2173.320 1095.160 2173.580 ;
        RECT 1095.360 2173.320 1095.620 2173.580 ;
        RECT 1096.740 2010.800 1097.000 2011.060 ;
        RECT 1313.860 2010.800 1314.120 2011.060 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3517.370 1095.100 3517.600 ;
        RECT 1094.500 3517.230 1095.100 3517.370 ;
        RECT 1094.500 3478.725 1094.640 3517.230 ;
        RECT 1094.430 3478.355 1094.710 3478.725 ;
        RECT 1096.270 3477.930 1096.550 3478.045 ;
        RECT 1095.880 3477.790 1096.550 3477.930 ;
        RECT 1095.880 3477.510 1096.020 3477.790 ;
        RECT 1096.270 3477.675 1096.550 3477.790 ;
        RECT 1095.820 3477.190 1096.080 3477.510 ;
        RECT 1095.360 3429.250 1095.620 3429.570 ;
        RECT 1095.420 3394.970 1095.560 3429.250 ;
        RECT 1094.960 3394.830 1095.560 3394.970 ;
        RECT 1094.960 3380.950 1095.100 3394.830 ;
        RECT 1094.900 3380.630 1095.160 3380.950 ;
        RECT 1095.360 3332.690 1095.620 3333.010 ;
        RECT 1095.420 3298.410 1095.560 3332.690 ;
        RECT 1095.420 3298.330 1096.020 3298.410 ;
        RECT 1095.420 3298.270 1096.080 3298.330 ;
        RECT 1095.820 3298.010 1096.080 3298.270 ;
        RECT 1096.740 3298.010 1097.000 3298.330 ;
        RECT 1096.800 3284.390 1096.940 3298.010 ;
        RECT 1096.740 3284.070 1097.000 3284.390 ;
        RECT 1096.280 3236.130 1096.540 3236.450 ;
        RECT 1096.340 3202.110 1096.480 3236.130 ;
        RECT 1096.280 3201.790 1096.540 3202.110 ;
        RECT 1095.360 3201.110 1095.620 3201.430 ;
        RECT 1095.420 3187.830 1095.560 3201.110 ;
        RECT 1095.360 3187.510 1095.620 3187.830 ;
        RECT 1095.820 3187.510 1096.080 3187.830 ;
        RECT 1095.880 3152.890 1096.020 3187.510 ;
        RECT 1095.880 3152.750 1096.940 3152.890 ;
        RECT 1096.800 3132.750 1096.940 3152.750 ;
        RECT 1096.740 3132.430 1097.000 3132.750 ;
        RECT 1096.740 3084.150 1097.000 3084.470 ;
        RECT 1096.800 3057.270 1096.940 3084.150 ;
        RECT 1096.740 3056.950 1097.000 3057.270 ;
        RECT 1095.360 3043.350 1095.620 3043.670 ;
        RECT 1095.420 3042.990 1095.560 3043.350 ;
        RECT 1095.360 3042.670 1095.620 3042.990 ;
        RECT 1096.280 3007.650 1096.540 3007.970 ;
        RECT 1096.340 2994.710 1096.480 3007.650 ;
        RECT 1096.280 2994.390 1096.540 2994.710 ;
        RECT 1095.820 2946.450 1096.080 2946.770 ;
        RECT 1095.880 2912.090 1096.020 2946.450 ;
        RECT 1094.900 2911.770 1095.160 2912.090 ;
        RECT 1095.820 2911.770 1096.080 2912.090 ;
        RECT 1094.960 2898.150 1095.100 2911.770 ;
        RECT 1094.900 2897.830 1095.160 2898.150 ;
        RECT 1094.440 2849.550 1094.700 2849.870 ;
        RECT 1094.500 2815.530 1094.640 2849.550 ;
        RECT 1094.440 2815.210 1094.700 2815.530 ;
        RECT 1094.900 2814.530 1095.160 2814.850 ;
        RECT 1094.960 2801.330 1095.100 2814.530 ;
        RECT 1094.500 2801.190 1095.100 2801.330 ;
        RECT 1094.500 2767.250 1094.640 2801.190 ;
        RECT 1094.440 2766.930 1094.700 2767.250 ;
        RECT 1094.440 2752.990 1094.700 2753.310 ;
        RECT 1094.500 2718.970 1094.640 2752.990 ;
        RECT 1094.440 2718.650 1094.700 2718.970 ;
        RECT 1094.900 2717.970 1095.160 2718.290 ;
        RECT 1094.960 2704.885 1095.100 2717.970 ;
        RECT 1094.890 2704.515 1095.170 2704.885 ;
        RECT 1095.810 2704.515 1096.090 2704.885 ;
        RECT 1095.880 2669.410 1096.020 2704.515 ;
        RECT 1094.960 2669.270 1096.020 2669.410 ;
        RECT 1094.960 2656.605 1095.100 2669.270 ;
        RECT 1094.890 2656.235 1095.170 2656.605 ;
        RECT 1095.810 2656.235 1096.090 2656.605 ;
        RECT 1095.880 2621.730 1096.020 2656.235 ;
        RECT 1094.900 2621.410 1095.160 2621.730 ;
        RECT 1095.820 2621.410 1096.080 2621.730 ;
        RECT 1094.960 2608.325 1095.100 2621.410 ;
        RECT 1093.970 2607.955 1094.250 2608.325 ;
        RECT 1094.890 2607.955 1095.170 2608.325 ;
        RECT 1094.040 2573.450 1094.180 2607.955 ;
        RECT 1093.980 2573.130 1094.240 2573.450 ;
        RECT 1095.360 2573.130 1095.620 2573.450 ;
        RECT 1095.420 2553.050 1095.560 2573.130 ;
        RECT 1095.360 2552.730 1095.620 2553.050 ;
        RECT 1095.360 2525.190 1095.620 2525.510 ;
        RECT 1095.420 2463.630 1095.560 2525.190 ;
        RECT 1095.360 2463.310 1095.620 2463.630 ;
        RECT 1095.820 2463.310 1096.080 2463.630 ;
        RECT 1095.880 2429.290 1096.020 2463.310 ;
        RECT 1095.820 2428.970 1096.080 2429.290 ;
        RECT 1096.280 2428.290 1096.540 2428.610 ;
        RECT 1096.340 2366.925 1096.480 2428.290 ;
        RECT 1094.890 2366.555 1095.170 2366.925 ;
        RECT 1096.270 2366.555 1096.550 2366.925 ;
        RECT 1094.960 2332.390 1095.100 2366.555 ;
        RECT 1094.900 2332.070 1095.160 2332.390 ;
        RECT 1096.740 2331.390 1097.000 2331.710 ;
        RECT 1096.800 2283.850 1096.940 2331.390 ;
        RECT 1095.420 2283.710 1096.940 2283.850 ;
        RECT 1095.420 2270.170 1095.560 2283.710 ;
        RECT 1095.360 2269.850 1095.620 2270.170 ;
        RECT 1094.900 2221.910 1095.160 2222.230 ;
        RECT 1094.960 2187.290 1095.100 2221.910 ;
        RECT 1094.960 2187.150 1095.560 2187.290 ;
        RECT 1095.420 2173.610 1095.560 2187.150 ;
        RECT 1094.900 2173.290 1095.160 2173.610 ;
        RECT 1095.360 2173.290 1095.620 2173.610 ;
        RECT 1094.960 2125.525 1095.100 2173.290 ;
        RECT 1094.890 2125.155 1095.170 2125.525 ;
        RECT 1096.730 2125.155 1097.010 2125.525 ;
        RECT 1096.800 2011.090 1096.940 2125.155 ;
        RECT 1096.740 2010.770 1097.000 2011.090 ;
        RECT 1313.860 2010.770 1314.120 2011.090 ;
        RECT 1313.920 2000.000 1314.060 2010.770 ;
        RECT 1313.760 1999.540 1314.060 2000.000 ;
        RECT 1313.760 1996.000 1314.040 1999.540 ;
      LAYER via2 ;
        RECT 1094.430 3478.400 1094.710 3478.680 ;
        RECT 1096.270 3477.720 1096.550 3478.000 ;
        RECT 1094.890 2704.560 1095.170 2704.840 ;
        RECT 1095.810 2704.560 1096.090 2704.840 ;
        RECT 1094.890 2656.280 1095.170 2656.560 ;
        RECT 1095.810 2656.280 1096.090 2656.560 ;
        RECT 1093.970 2608.000 1094.250 2608.280 ;
        RECT 1094.890 2608.000 1095.170 2608.280 ;
        RECT 1094.890 2366.600 1095.170 2366.880 ;
        RECT 1096.270 2366.600 1096.550 2366.880 ;
        RECT 1094.890 2125.200 1095.170 2125.480 ;
        RECT 1096.730 2125.200 1097.010 2125.480 ;
      LAYER met3 ;
        RECT 1094.405 3478.690 1094.735 3478.705 ;
        RECT 1094.405 3478.390 1097.250 3478.690 ;
        RECT 1094.405 3478.375 1094.735 3478.390 ;
        RECT 1096.245 3478.010 1096.575 3478.025 ;
        RECT 1096.950 3478.010 1097.250 3478.390 ;
        RECT 1096.245 3477.710 1097.250 3478.010 ;
        RECT 1096.245 3477.695 1096.575 3477.710 ;
        RECT 1094.865 2704.850 1095.195 2704.865 ;
        RECT 1095.785 2704.850 1096.115 2704.865 ;
        RECT 1094.865 2704.550 1096.115 2704.850 ;
        RECT 1094.865 2704.535 1095.195 2704.550 ;
        RECT 1095.785 2704.535 1096.115 2704.550 ;
        RECT 1094.865 2656.570 1095.195 2656.585 ;
        RECT 1095.785 2656.570 1096.115 2656.585 ;
        RECT 1094.865 2656.270 1096.115 2656.570 ;
        RECT 1094.865 2656.255 1095.195 2656.270 ;
        RECT 1095.785 2656.255 1096.115 2656.270 ;
        RECT 1093.945 2608.290 1094.275 2608.305 ;
        RECT 1094.865 2608.290 1095.195 2608.305 ;
        RECT 1093.945 2607.990 1095.195 2608.290 ;
        RECT 1093.945 2607.975 1094.275 2607.990 ;
        RECT 1094.865 2607.975 1095.195 2607.990 ;
        RECT 1094.865 2366.890 1095.195 2366.905 ;
        RECT 1096.245 2366.890 1096.575 2366.905 ;
        RECT 1094.865 2366.590 1096.575 2366.890 ;
        RECT 1094.865 2366.575 1095.195 2366.590 ;
        RECT 1096.245 2366.575 1096.575 2366.590 ;
        RECT 1094.865 2125.490 1095.195 2125.505 ;
        RECT 1096.705 2125.490 1097.035 2125.505 ;
        RECT 1094.865 2125.190 1097.035 2125.490 ;
        RECT 1094.865 2125.175 1095.195 2125.190 ;
        RECT 1096.705 2125.175 1097.035 2125.190 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 771.565 3381.045 771.735 3429.155 ;
        RECT 771.565 2898.585 771.735 2946.355 ;
        RECT 772.025 2608.225 772.195 2656.335 ;
        RECT 772.025 2511.665 772.195 2559.775 ;
        RECT 771.105 2221.985 771.275 2270.095 ;
        RECT 772.025 2138.685 772.195 2173.535 ;
        RECT 771.565 2028.525 771.735 2076.975 ;
      LAYER mcon ;
        RECT 771.565 3428.985 771.735 3429.155 ;
        RECT 771.565 2946.185 771.735 2946.355 ;
        RECT 772.025 2656.165 772.195 2656.335 ;
        RECT 772.025 2559.605 772.195 2559.775 ;
        RECT 771.105 2269.925 771.275 2270.095 ;
        RECT 772.025 2173.365 772.195 2173.535 ;
        RECT 771.565 2076.805 771.735 2076.975 ;
      LAYER met1 ;
        RECT 770.570 3477.760 770.890 3477.820 ;
        RECT 771.030 3477.760 771.350 3477.820 ;
        RECT 770.570 3477.620 771.350 3477.760 ;
        RECT 770.570 3477.560 770.890 3477.620 ;
        RECT 771.030 3477.560 771.350 3477.620 ;
        RECT 771.030 3443.080 771.350 3443.140 ;
        RECT 771.950 3443.080 772.270 3443.140 ;
        RECT 771.030 3442.940 772.270 3443.080 ;
        RECT 771.030 3442.880 771.350 3442.940 ;
        RECT 771.950 3442.880 772.270 3442.940 ;
        RECT 771.505 3429.140 771.795 3429.185 ;
        RECT 771.950 3429.140 772.270 3429.200 ;
        RECT 771.505 3429.000 772.270 3429.140 ;
        RECT 771.505 3428.955 771.795 3429.000 ;
        RECT 771.950 3428.940 772.270 3429.000 ;
        RECT 771.490 3381.200 771.810 3381.260 ;
        RECT 771.295 3381.060 771.810 3381.200 ;
        RECT 771.490 3381.000 771.810 3381.060 ;
        RECT 771.490 3367.600 771.810 3367.660 ;
        RECT 772.410 3367.600 772.730 3367.660 ;
        RECT 771.490 3367.460 772.730 3367.600 ;
        RECT 771.490 3367.400 771.810 3367.460 ;
        RECT 772.410 3367.400 772.730 3367.460 ;
        RECT 771.490 3270.700 771.810 3270.760 ;
        RECT 772.410 3270.700 772.730 3270.760 ;
        RECT 771.490 3270.560 772.730 3270.700 ;
        RECT 771.490 3270.500 771.810 3270.560 ;
        RECT 772.410 3270.500 772.730 3270.560 ;
        RECT 771.490 3174.140 771.810 3174.200 ;
        RECT 772.410 3174.140 772.730 3174.200 ;
        RECT 771.490 3174.000 772.730 3174.140 ;
        RECT 771.490 3173.940 771.810 3174.000 ;
        RECT 772.410 3173.940 772.730 3174.000 ;
        RECT 771.490 3077.580 771.810 3077.640 ;
        RECT 772.410 3077.580 772.730 3077.640 ;
        RECT 771.490 3077.440 772.730 3077.580 ;
        RECT 771.490 3077.380 771.810 3077.440 ;
        RECT 772.410 3077.380 772.730 3077.440 ;
        RECT 771.490 2981.020 771.810 2981.080 ;
        RECT 772.410 2981.020 772.730 2981.080 ;
        RECT 771.490 2980.880 772.730 2981.020 ;
        RECT 771.490 2980.820 771.810 2980.880 ;
        RECT 772.410 2980.820 772.730 2980.880 ;
        RECT 771.490 2946.340 771.810 2946.400 ;
        RECT 771.295 2946.200 771.810 2946.340 ;
        RECT 771.490 2946.140 771.810 2946.200 ;
        RECT 771.490 2898.740 771.810 2898.800 ;
        RECT 771.295 2898.600 771.810 2898.740 ;
        RECT 771.490 2898.540 771.810 2898.600 ;
        RECT 771.030 2898.060 771.350 2898.120 ;
        RECT 771.950 2898.060 772.270 2898.120 ;
        RECT 771.030 2897.920 772.270 2898.060 ;
        RECT 771.030 2897.860 771.350 2897.920 ;
        RECT 771.950 2897.860 772.270 2897.920 ;
        RECT 771.030 2814.760 771.350 2814.820 ;
        RECT 771.950 2814.760 772.270 2814.820 ;
        RECT 771.030 2814.620 772.270 2814.760 ;
        RECT 771.030 2814.560 771.350 2814.620 ;
        RECT 771.950 2814.560 772.270 2814.620 ;
        RECT 771.950 2656.320 772.270 2656.380 ;
        RECT 771.755 2656.180 772.270 2656.320 ;
        RECT 771.950 2656.120 772.270 2656.180 ;
        RECT 771.965 2608.380 772.255 2608.425 ;
        RECT 772.410 2608.380 772.730 2608.440 ;
        RECT 771.965 2608.240 772.730 2608.380 ;
        RECT 771.965 2608.195 772.255 2608.240 ;
        RECT 772.410 2608.180 772.730 2608.240 ;
        RECT 771.950 2559.760 772.270 2559.820 ;
        RECT 771.755 2559.620 772.270 2559.760 ;
        RECT 771.950 2559.560 772.270 2559.620 ;
        RECT 771.965 2511.820 772.255 2511.865 ;
        RECT 772.410 2511.820 772.730 2511.880 ;
        RECT 771.965 2511.680 772.730 2511.820 ;
        RECT 771.965 2511.635 772.255 2511.680 ;
        RECT 772.410 2511.620 772.730 2511.680 ;
        RECT 771.030 2463.200 771.350 2463.260 ;
        RECT 771.950 2463.200 772.270 2463.260 ;
        RECT 771.030 2463.060 772.270 2463.200 ;
        RECT 771.030 2463.000 771.350 2463.060 ;
        RECT 771.950 2463.000 772.270 2463.060 ;
        RECT 771.490 2332.300 771.810 2332.360 ;
        RECT 772.410 2332.300 772.730 2332.360 ;
        RECT 771.490 2332.160 772.730 2332.300 ;
        RECT 771.490 2332.100 771.810 2332.160 ;
        RECT 772.410 2332.100 772.730 2332.160 ;
        RECT 771.045 2270.080 771.335 2270.125 ;
        RECT 771.490 2270.080 771.810 2270.140 ;
        RECT 771.045 2269.940 771.810 2270.080 ;
        RECT 771.045 2269.895 771.335 2269.940 ;
        RECT 771.490 2269.880 771.810 2269.940 ;
        RECT 771.030 2222.140 771.350 2222.200 ;
        RECT 770.835 2222.000 771.350 2222.140 ;
        RECT 771.030 2221.940 771.350 2222.000 ;
        RECT 771.950 2173.520 772.270 2173.580 ;
        RECT 771.755 2173.380 772.270 2173.520 ;
        RECT 771.950 2173.320 772.270 2173.380 ;
        RECT 771.950 2138.840 772.270 2138.900 ;
        RECT 771.755 2138.700 772.270 2138.840 ;
        RECT 771.950 2138.640 772.270 2138.700 ;
        RECT 771.490 2076.960 771.810 2077.020 ;
        RECT 771.295 2076.820 771.810 2076.960 ;
        RECT 771.490 2076.760 771.810 2076.820 ;
        RECT 771.505 2028.680 771.795 2028.725 ;
        RECT 771.950 2028.680 772.270 2028.740 ;
        RECT 771.505 2028.540 772.270 2028.680 ;
        RECT 771.505 2028.495 771.795 2028.540 ;
        RECT 771.950 2028.480 772.270 2028.540 ;
        RECT 771.950 2014.400 772.270 2014.460 ;
        RECT 1321.650 2014.400 1321.970 2014.460 ;
        RECT 771.950 2014.260 1321.970 2014.400 ;
        RECT 771.950 2014.200 772.270 2014.260 ;
        RECT 1321.650 2014.200 1321.970 2014.260 ;
      LAYER via ;
        RECT 770.600 3477.560 770.860 3477.820 ;
        RECT 771.060 3477.560 771.320 3477.820 ;
        RECT 771.060 3442.880 771.320 3443.140 ;
        RECT 771.980 3442.880 772.240 3443.140 ;
        RECT 771.980 3428.940 772.240 3429.200 ;
        RECT 771.520 3381.000 771.780 3381.260 ;
        RECT 771.520 3367.400 771.780 3367.660 ;
        RECT 772.440 3367.400 772.700 3367.660 ;
        RECT 771.520 3270.500 771.780 3270.760 ;
        RECT 772.440 3270.500 772.700 3270.760 ;
        RECT 771.520 3173.940 771.780 3174.200 ;
        RECT 772.440 3173.940 772.700 3174.200 ;
        RECT 771.520 3077.380 771.780 3077.640 ;
        RECT 772.440 3077.380 772.700 3077.640 ;
        RECT 771.520 2980.820 771.780 2981.080 ;
        RECT 772.440 2980.820 772.700 2981.080 ;
        RECT 771.520 2946.140 771.780 2946.400 ;
        RECT 771.520 2898.540 771.780 2898.800 ;
        RECT 771.060 2897.860 771.320 2898.120 ;
        RECT 771.980 2897.860 772.240 2898.120 ;
        RECT 771.060 2814.560 771.320 2814.820 ;
        RECT 771.980 2814.560 772.240 2814.820 ;
        RECT 771.980 2656.120 772.240 2656.380 ;
        RECT 772.440 2608.180 772.700 2608.440 ;
        RECT 771.980 2559.560 772.240 2559.820 ;
        RECT 772.440 2511.620 772.700 2511.880 ;
        RECT 771.060 2463.000 771.320 2463.260 ;
        RECT 771.980 2463.000 772.240 2463.260 ;
        RECT 771.520 2332.100 771.780 2332.360 ;
        RECT 772.440 2332.100 772.700 2332.360 ;
        RECT 771.520 2269.880 771.780 2270.140 ;
        RECT 771.060 2221.940 771.320 2222.200 ;
        RECT 771.980 2173.320 772.240 2173.580 ;
        RECT 771.980 2138.640 772.240 2138.900 ;
        RECT 771.520 2076.760 771.780 2077.020 ;
        RECT 771.980 2028.480 772.240 2028.740 ;
        RECT 771.980 2014.200 772.240 2014.460 ;
        RECT 1321.680 2014.200 1321.940 2014.460 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3477.850 770.800 3517.600 ;
        RECT 770.600 3477.530 770.860 3477.850 ;
        RECT 771.060 3477.530 771.320 3477.850 ;
        RECT 771.120 3443.170 771.260 3477.530 ;
        RECT 771.060 3442.850 771.320 3443.170 ;
        RECT 771.980 3442.850 772.240 3443.170 ;
        RECT 772.040 3429.230 772.180 3442.850 ;
        RECT 771.980 3428.910 772.240 3429.230 ;
        RECT 771.520 3380.970 771.780 3381.290 ;
        RECT 771.580 3367.690 771.720 3380.970 ;
        RECT 771.520 3367.370 771.780 3367.690 ;
        RECT 772.440 3367.370 772.700 3367.690 ;
        RECT 772.500 3318.810 772.640 3367.370 ;
        RECT 771.580 3318.670 772.640 3318.810 ;
        RECT 771.580 3270.790 771.720 3318.670 ;
        RECT 771.520 3270.470 771.780 3270.790 ;
        RECT 772.440 3270.470 772.700 3270.790 ;
        RECT 772.500 3222.250 772.640 3270.470 ;
        RECT 771.580 3222.110 772.640 3222.250 ;
        RECT 771.580 3174.230 771.720 3222.110 ;
        RECT 771.520 3173.910 771.780 3174.230 ;
        RECT 772.440 3173.910 772.700 3174.230 ;
        RECT 772.500 3125.690 772.640 3173.910 ;
        RECT 771.580 3125.550 772.640 3125.690 ;
        RECT 771.580 3077.670 771.720 3125.550 ;
        RECT 771.520 3077.350 771.780 3077.670 ;
        RECT 772.440 3077.350 772.700 3077.670 ;
        RECT 772.500 3029.130 772.640 3077.350 ;
        RECT 771.580 3028.990 772.640 3029.130 ;
        RECT 771.580 2981.110 771.720 3028.990 ;
        RECT 771.520 2980.790 771.780 2981.110 ;
        RECT 772.440 2980.850 772.700 2981.110 ;
        RECT 772.040 2980.790 772.700 2980.850 ;
        RECT 772.040 2980.710 772.640 2980.790 ;
        RECT 772.040 2959.770 772.180 2980.710 ;
        RECT 771.580 2959.630 772.180 2959.770 ;
        RECT 771.580 2946.430 771.720 2959.630 ;
        RECT 771.520 2946.110 771.780 2946.430 ;
        RECT 771.520 2898.570 771.780 2898.830 ;
        RECT 771.120 2898.510 771.780 2898.570 ;
        RECT 771.120 2898.430 771.720 2898.510 ;
        RECT 771.120 2898.150 771.260 2898.430 ;
        RECT 771.060 2897.830 771.320 2898.150 ;
        RECT 771.980 2897.830 772.240 2898.150 ;
        RECT 772.040 2814.850 772.180 2897.830 ;
        RECT 771.060 2814.530 771.320 2814.850 ;
        RECT 771.980 2814.530 772.240 2814.850 ;
        RECT 771.120 2766.650 771.260 2814.530 ;
        RECT 771.120 2766.510 771.720 2766.650 ;
        RECT 771.580 2719.050 771.720 2766.510 ;
        RECT 771.580 2718.910 772.640 2719.050 ;
        RECT 772.500 2670.090 772.640 2718.910 ;
        RECT 772.040 2669.950 772.640 2670.090 ;
        RECT 772.040 2656.410 772.180 2669.950 ;
        RECT 771.980 2656.090 772.240 2656.410 ;
        RECT 772.440 2608.150 772.700 2608.470 ;
        RECT 772.500 2573.530 772.640 2608.150 ;
        RECT 772.040 2573.390 772.640 2573.530 ;
        RECT 772.040 2559.850 772.180 2573.390 ;
        RECT 771.980 2559.530 772.240 2559.850 ;
        RECT 772.440 2511.590 772.700 2511.910 ;
        RECT 772.500 2476.970 772.640 2511.590 ;
        RECT 772.040 2476.830 772.640 2476.970 ;
        RECT 772.040 2463.290 772.180 2476.830 ;
        RECT 771.060 2462.970 771.320 2463.290 ;
        RECT 771.980 2462.970 772.240 2463.290 ;
        RECT 771.120 2415.205 771.260 2462.970 ;
        RECT 771.050 2414.835 771.330 2415.205 ;
        RECT 772.430 2414.835 772.710 2415.205 ;
        RECT 772.500 2380.410 772.640 2414.835 ;
        RECT 771.580 2380.270 772.640 2380.410 ;
        RECT 771.580 2332.390 771.720 2380.270 ;
        RECT 771.520 2332.070 771.780 2332.390 ;
        RECT 772.440 2332.070 772.700 2332.390 ;
        RECT 772.500 2283.850 772.640 2332.070 ;
        RECT 771.580 2283.710 772.640 2283.850 ;
        RECT 771.580 2270.170 771.720 2283.710 ;
        RECT 771.520 2269.850 771.780 2270.170 ;
        RECT 771.060 2221.910 771.320 2222.230 ;
        RECT 771.120 2187.290 771.260 2221.910 ;
        RECT 771.120 2187.150 772.180 2187.290 ;
        RECT 772.040 2173.610 772.180 2187.150 ;
        RECT 771.980 2173.290 772.240 2173.610 ;
        RECT 771.980 2138.610 772.240 2138.930 ;
        RECT 772.040 2125.410 772.180 2138.610 ;
        RECT 772.040 2125.270 772.640 2125.410 ;
        RECT 772.500 2090.730 772.640 2125.270 ;
        RECT 771.580 2090.590 772.640 2090.730 ;
        RECT 771.580 2077.050 771.720 2090.590 ;
        RECT 771.520 2076.730 771.780 2077.050 ;
        RECT 771.980 2028.450 772.240 2028.770 ;
        RECT 772.040 2014.490 772.180 2028.450 ;
        RECT 771.980 2014.170 772.240 2014.490 ;
        RECT 1321.680 2014.170 1321.940 2014.490 ;
        RECT 1321.740 2000.000 1321.880 2014.170 ;
        RECT 1321.580 1999.540 1321.880 2000.000 ;
        RECT 1321.580 1996.000 1321.860 1999.540 ;
      LAYER via2 ;
        RECT 771.050 2414.880 771.330 2415.160 ;
        RECT 772.430 2414.880 772.710 2415.160 ;
      LAYER met3 ;
        RECT 771.025 2415.170 771.355 2415.185 ;
        RECT 772.405 2415.170 772.735 2415.185 ;
        RECT 771.025 2414.870 772.735 2415.170 ;
        RECT 771.025 2414.855 771.355 2414.870 ;
        RECT 772.405 2414.855 772.735 2414.870 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3498.500 446.130 3498.560 ;
        RECT 448.110 3498.500 448.430 3498.560 ;
        RECT 445.810 3498.360 448.430 3498.500 ;
        RECT 445.810 3498.300 446.130 3498.360 ;
        RECT 448.110 3498.300 448.430 3498.360 ;
        RECT 448.110 2013.720 448.430 2013.780 ;
        RECT 448.110 2013.580 1291.520 2013.720 ;
        RECT 448.110 2013.520 448.430 2013.580 ;
        RECT 1291.380 2013.380 1291.520 2013.580 ;
        RECT 1329.470 2013.380 1329.790 2013.440 ;
        RECT 1291.380 2013.240 1329.790 2013.380 ;
        RECT 1329.470 2013.180 1329.790 2013.240 ;
      LAYER via ;
        RECT 445.840 3498.300 446.100 3498.560 ;
        RECT 448.140 3498.300 448.400 3498.560 ;
        RECT 448.140 2013.520 448.400 2013.780 ;
        RECT 1329.500 2013.180 1329.760 2013.440 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3498.590 446.040 3517.600 ;
        RECT 445.840 3498.270 446.100 3498.590 ;
        RECT 448.140 3498.270 448.400 3498.590 ;
        RECT 448.200 2013.810 448.340 3498.270 ;
        RECT 448.140 2013.490 448.400 2013.810 ;
        RECT 1329.500 2013.150 1329.760 2013.470 ;
        RECT 1329.560 2000.000 1329.700 2013.150 ;
        RECT 1329.400 1999.540 1329.700 2000.000 ;
        RECT 1329.400 1996.000 1329.680 1999.540 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 123.810 2013.040 124.130 2013.100 ;
        RECT 1290.370 2013.040 1290.690 2013.100 ;
        RECT 123.810 2012.900 1290.690 2013.040 ;
        RECT 123.810 2012.840 124.130 2012.900 ;
        RECT 1290.370 2012.840 1290.690 2012.900 ;
        RECT 1337.750 2012.700 1338.070 2012.760 ;
        RECT 1314.380 2012.560 1338.070 2012.700 ;
        RECT 1306.010 2012.360 1306.330 2012.420 ;
        RECT 1314.380 2012.360 1314.520 2012.560 ;
        RECT 1337.750 2012.500 1338.070 2012.560 ;
        RECT 1306.010 2012.220 1314.520 2012.360 ;
        RECT 1306.010 2012.160 1306.330 2012.220 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 123.840 2012.840 124.100 2013.100 ;
        RECT 1290.400 2012.840 1290.660 2013.100 ;
        RECT 1306.040 2012.160 1306.300 2012.420 ;
        RECT 1337.780 2012.500 1338.040 2012.760 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 2013.130 124.040 3498.270 ;
        RECT 123.840 2012.810 124.100 2013.130 ;
        RECT 1290.400 2012.810 1290.660 2013.130 ;
        RECT 1290.460 2012.645 1290.600 2012.810 ;
        RECT 1290.390 2012.275 1290.670 2012.645 ;
        RECT 1306.030 2012.275 1306.310 2012.645 ;
        RECT 1337.780 2012.470 1338.040 2012.790 ;
        RECT 1306.040 2012.130 1306.300 2012.275 ;
        RECT 1337.840 2000.000 1337.980 2012.470 ;
        RECT 1337.680 1999.540 1337.980 2000.000 ;
        RECT 1337.680 1996.000 1337.960 1999.540 ;
      LAYER via2 ;
        RECT 1290.390 2012.320 1290.670 2012.600 ;
        RECT 1306.030 2012.320 1306.310 2012.600 ;
      LAYER met3 ;
        RECT 1290.365 2012.610 1290.695 2012.625 ;
        RECT 1306.005 2012.610 1306.335 2012.625 ;
        RECT 1290.365 2012.310 1306.335 2012.610 ;
        RECT 1290.365 2012.295 1290.695 2012.310 ;
        RECT 1306.005 2012.295 1306.335 2012.310 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 3339.720 17.870 3339.780 ;
        RECT 1314.290 3339.720 1314.610 3339.780 ;
        RECT 17.550 3339.580 1314.610 3339.720 ;
        RECT 17.550 3339.520 17.870 3339.580 ;
        RECT 1314.290 3339.520 1314.610 3339.580 ;
        RECT 1314.750 2012.360 1315.070 2012.420 ;
        RECT 1345.570 2012.360 1345.890 2012.420 ;
        RECT 1314.750 2012.220 1345.890 2012.360 ;
        RECT 1314.750 2012.160 1315.070 2012.220 ;
        RECT 1345.570 2012.160 1345.890 2012.220 ;
      LAYER via ;
        RECT 17.580 3339.520 17.840 3339.780 ;
        RECT 1314.320 3339.520 1314.580 3339.780 ;
        RECT 1314.780 2012.160 1315.040 2012.420 ;
        RECT 1345.600 2012.160 1345.860 2012.420 ;
      LAYER met2 ;
        RECT 17.570 3339.635 17.850 3340.005 ;
        RECT 17.580 3339.490 17.840 3339.635 ;
        RECT 1314.320 3339.490 1314.580 3339.810 ;
        RECT 1314.380 2013.890 1314.520 3339.490 ;
        RECT 1314.380 2013.750 1314.980 2013.890 ;
        RECT 1314.840 2012.450 1314.980 2013.750 ;
        RECT 1314.780 2012.130 1315.040 2012.450 ;
        RECT 1345.600 2012.130 1345.860 2012.450 ;
        RECT 1345.660 2000.000 1345.800 2012.130 ;
        RECT 1345.500 1999.540 1345.800 2000.000 ;
        RECT 1345.500 1996.000 1345.780 1999.540 ;
      LAYER via2 ;
        RECT 17.570 3339.680 17.850 3339.960 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.545 3339.970 17.875 3339.985 ;
        RECT -4.800 3339.670 17.875 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.545 3339.655 17.875 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 3050.040 18.330 3050.100 ;
        RECT 1321.190 3050.040 1321.510 3050.100 ;
        RECT 18.010 3049.900 1321.510 3050.040 ;
        RECT 18.010 3049.840 18.330 3049.900 ;
        RECT 1321.190 3049.840 1321.510 3049.900 ;
        RECT 1321.190 2014.060 1321.510 2014.120 ;
        RECT 1353.390 2014.060 1353.710 2014.120 ;
        RECT 1321.190 2013.920 1353.710 2014.060 ;
        RECT 1321.190 2013.860 1321.510 2013.920 ;
        RECT 1353.390 2013.860 1353.710 2013.920 ;
      LAYER via ;
        RECT 18.040 3049.840 18.300 3050.100 ;
        RECT 1321.220 3049.840 1321.480 3050.100 ;
        RECT 1321.220 2013.860 1321.480 2014.120 ;
        RECT 1353.420 2013.860 1353.680 2014.120 ;
      LAYER met2 ;
        RECT 18.030 3051.995 18.310 3052.365 ;
        RECT 18.100 3050.130 18.240 3051.995 ;
        RECT 18.040 3049.810 18.300 3050.130 ;
        RECT 1321.220 3049.810 1321.480 3050.130 ;
        RECT 1321.280 2014.150 1321.420 3049.810 ;
        RECT 1321.220 2013.830 1321.480 2014.150 ;
        RECT 1353.420 2013.830 1353.680 2014.150 ;
        RECT 1353.480 2000.000 1353.620 2013.830 ;
        RECT 1353.320 1999.540 1353.620 2000.000 ;
        RECT 1353.320 1996.000 1353.600 1999.540 ;
      LAYER via2 ;
        RECT 18.030 3052.040 18.310 3052.320 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 18.005 3052.330 18.335 3052.345 ;
        RECT -4.800 3052.030 18.335 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 18.005 3052.015 18.335 3052.030 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2760.360 16.950 2760.420 ;
        RECT 1328.090 2760.360 1328.410 2760.420 ;
        RECT 16.630 2760.220 1328.410 2760.360 ;
        RECT 16.630 2760.160 16.950 2760.220 ;
        RECT 1328.090 2760.160 1328.410 2760.220 ;
        RECT 1328.090 2013.720 1328.410 2013.780 ;
        RECT 1361.210 2013.720 1361.530 2013.780 ;
        RECT 1328.090 2013.580 1361.530 2013.720 ;
        RECT 1328.090 2013.520 1328.410 2013.580 ;
        RECT 1361.210 2013.520 1361.530 2013.580 ;
      LAYER via ;
        RECT 16.660 2760.160 16.920 2760.420 ;
        RECT 1328.120 2760.160 1328.380 2760.420 ;
        RECT 1328.120 2013.520 1328.380 2013.780 ;
        RECT 1361.240 2013.520 1361.500 2013.780 ;
      LAYER met2 ;
        RECT 16.650 2765.035 16.930 2765.405 ;
        RECT 16.720 2760.450 16.860 2765.035 ;
        RECT 16.660 2760.130 16.920 2760.450 ;
        RECT 1328.120 2760.130 1328.380 2760.450 ;
        RECT 1328.180 2013.810 1328.320 2760.130 ;
        RECT 1328.120 2013.490 1328.380 2013.810 ;
        RECT 1361.240 2013.490 1361.500 2013.810 ;
        RECT 1361.300 2000.000 1361.440 2013.490 ;
        RECT 1361.140 1999.540 1361.440 2000.000 ;
        RECT 1361.140 1996.000 1361.420 1999.540 ;
      LAYER via2 ;
        RECT 16.650 2765.080 16.930 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 16.625 2765.370 16.955 2765.385 ;
        RECT -4.800 2765.070 16.955 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 16.625 2765.055 16.955 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2477.480 16.950 2477.540 ;
        RECT 1334.990 2477.480 1335.310 2477.540 ;
        RECT 16.630 2477.340 1335.310 2477.480 ;
        RECT 16.630 2477.280 16.950 2477.340 ;
        RECT 1334.990 2477.280 1335.310 2477.340 ;
        RECT 1334.990 2013.040 1335.310 2013.100 ;
        RECT 1369.030 2013.040 1369.350 2013.100 ;
        RECT 1334.990 2012.900 1369.350 2013.040 ;
        RECT 1334.990 2012.840 1335.310 2012.900 ;
        RECT 1369.030 2012.840 1369.350 2012.900 ;
      LAYER via ;
        RECT 16.660 2477.280 16.920 2477.540 ;
        RECT 1335.020 2477.280 1335.280 2477.540 ;
        RECT 1335.020 2012.840 1335.280 2013.100 ;
        RECT 1369.060 2012.840 1369.320 2013.100 ;
      LAYER met2 ;
        RECT 16.650 2477.395 16.930 2477.765 ;
        RECT 16.660 2477.250 16.920 2477.395 ;
        RECT 1335.020 2477.250 1335.280 2477.570 ;
        RECT 1335.080 2013.130 1335.220 2477.250 ;
        RECT 1335.020 2012.810 1335.280 2013.130 ;
        RECT 1369.060 2012.810 1369.320 2013.130 ;
        RECT 1369.120 2000.000 1369.260 2012.810 ;
        RECT 1368.960 1999.540 1369.260 2000.000 ;
        RECT 1368.960 1996.000 1369.240 1999.540 ;
      LAYER via2 ;
        RECT 16.650 2477.440 16.930 2477.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 16.625 2477.730 16.955 2477.745 ;
        RECT -4.800 2477.430 16.955 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 16.625 2477.415 16.955 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2187.460 16.950 2187.520 ;
        RECT 1348.790 2187.460 1349.110 2187.520 ;
        RECT 16.630 2187.320 1349.110 2187.460 ;
        RECT 16.630 2187.260 16.950 2187.320 ;
        RECT 1348.790 2187.260 1349.110 2187.320 ;
        RECT 1348.790 2011.000 1349.110 2011.060 ;
        RECT 1376.850 2011.000 1377.170 2011.060 ;
        RECT 1348.790 2010.860 1377.170 2011.000 ;
        RECT 1348.790 2010.800 1349.110 2010.860 ;
        RECT 1376.850 2010.800 1377.170 2010.860 ;
      LAYER via ;
        RECT 16.660 2187.260 16.920 2187.520 ;
        RECT 1348.820 2187.260 1349.080 2187.520 ;
        RECT 1348.820 2010.800 1349.080 2011.060 ;
        RECT 1376.880 2010.800 1377.140 2011.060 ;
      LAYER met2 ;
        RECT 16.650 2189.755 16.930 2190.125 ;
        RECT 16.720 2187.550 16.860 2189.755 ;
        RECT 16.660 2187.230 16.920 2187.550 ;
        RECT 1348.820 2187.230 1349.080 2187.550 ;
        RECT 1348.880 2011.090 1349.020 2187.230 ;
        RECT 1348.820 2010.770 1349.080 2011.090 ;
        RECT 1376.880 2010.770 1377.140 2011.090 ;
        RECT 1376.940 2000.000 1377.080 2010.770 ;
        RECT 1376.780 1999.540 1377.080 2000.000 ;
        RECT 1376.780 1996.000 1377.060 1999.540 ;
      LAYER via2 ;
        RECT 16.650 2189.800 16.930 2190.080 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 16.625 2190.090 16.955 2190.105 ;
        RECT -4.800 2189.790 16.955 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 16.625 2189.775 16.955 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1904.240 17.410 1904.300 ;
        RECT 1128.450 1904.240 1128.770 1904.300 ;
        RECT 17.090 1904.100 1128.770 1904.240 ;
        RECT 17.090 1904.040 17.410 1904.100 ;
        RECT 1128.450 1904.040 1128.770 1904.100 ;
      LAYER via ;
        RECT 17.120 1904.040 17.380 1904.300 ;
        RECT 1128.480 1904.040 1128.740 1904.300 ;
      LAYER met2 ;
        RECT 1384.230 1996.890 1384.510 1997.005 ;
        RECT 1385.060 1996.890 1385.340 2000.000 ;
        RECT 1384.230 1996.750 1385.340 1996.890 ;
        RECT 1384.230 1996.635 1384.510 1996.750 ;
        RECT 1385.060 1996.000 1385.340 1996.750 ;
        RECT 1128.470 1993.235 1128.750 1993.605 ;
        RECT 1128.540 1904.330 1128.680 1993.235 ;
        RECT 17.120 1904.010 17.380 1904.330 ;
        RECT 1128.480 1904.010 1128.740 1904.330 ;
        RECT 17.180 1903.165 17.320 1904.010 ;
        RECT 17.110 1902.795 17.390 1903.165 ;
      LAYER via2 ;
        RECT 1384.230 1996.680 1384.510 1996.960 ;
        RECT 1128.470 1993.280 1128.750 1993.560 ;
        RECT 17.110 1902.840 17.390 1903.120 ;
      LAYER met3 ;
        RECT 1384.205 1996.980 1384.535 1996.985 ;
        RECT 1383.950 1996.970 1384.535 1996.980 ;
        RECT 1383.750 1996.670 1384.535 1996.970 ;
        RECT 1383.950 1996.660 1384.535 1996.670 ;
        RECT 1384.205 1996.655 1384.535 1996.660 ;
        RECT 1128.445 1993.570 1128.775 1993.585 ;
        RECT 1383.950 1993.570 1384.330 1993.580 ;
        RECT 1128.445 1993.270 1384.330 1993.570 ;
        RECT 1128.445 1993.255 1128.775 1993.270 ;
        RECT 1383.950 1993.260 1384.330 1993.270 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 17.085 1903.130 17.415 1903.145 ;
        RECT -4.800 1902.830 17.415 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 17.085 1902.815 17.415 1902.830 ;
      LAYER via3 ;
        RECT 1383.980 1996.660 1384.300 1996.980 ;
        RECT 1383.980 1993.260 1384.300 1993.580 ;
      LAYER met4 ;
        RECT 1383.975 1996.655 1384.305 1996.985 ;
        RECT 1383.990 1993.585 1384.290 1996.655 ;
        RECT 1383.975 1993.255 1384.305 1993.585 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1172.685 1995.205 1172.855 1996.395 ;
      LAYER mcon ;
        RECT 1172.685 1996.225 1172.855 1996.395 ;
      LAYER met1 ;
        RECT 1172.610 1996.380 1172.930 1996.440 ;
        RECT 1172.415 1996.240 1172.930 1996.380 ;
        RECT 1172.610 1996.180 1172.930 1996.240 ;
        RECT 1172.625 1995.360 1172.915 1995.405 ;
        RECT 1562.690 1995.360 1563.010 1995.420 ;
        RECT 1172.625 1995.220 1563.010 1995.360 ;
        RECT 1172.625 1995.175 1172.915 1995.220 ;
        RECT 1562.690 1995.160 1563.010 1995.220 ;
        RECT 1562.690 620.740 1563.010 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 1562.690 620.600 2901.150 620.740 ;
        RECT 1562.690 620.540 1563.010 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 1172.640 1996.180 1172.900 1996.440 ;
        RECT 1562.720 1995.160 1562.980 1995.420 ;
        RECT 1562.720 620.540 1562.980 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 1171.620 1996.890 1171.900 2000.000 ;
        RECT 1171.620 1996.750 1172.840 1996.890 ;
        RECT 1171.620 1996.000 1171.900 1996.750 ;
        RECT 1172.700 1996.470 1172.840 1996.750 ;
        RECT 1172.640 1996.150 1172.900 1996.470 ;
        RECT 1562.720 1995.130 1562.980 1995.450 ;
        RECT 1562.780 620.830 1562.920 1995.130 ;
        RECT 1562.720 620.510 1562.980 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1240.765 2008.805 1241.855 2008.975 ;
      LAYER mcon ;
        RECT 1241.685 2008.805 1241.855 2008.975 ;
      LAYER met1 ;
        RECT 19.850 2008.960 20.170 2009.020 ;
        RECT 1240.705 2008.960 1240.995 2009.005 ;
        RECT 19.850 2008.820 1240.995 2008.960 ;
        RECT 19.850 2008.760 20.170 2008.820 ;
        RECT 1240.705 2008.775 1240.995 2008.820 ;
        RECT 1241.625 2008.960 1241.915 2009.005 ;
        RECT 1392.950 2008.960 1393.270 2009.020 ;
        RECT 1241.625 2008.820 1393.270 2008.960 ;
        RECT 1241.625 2008.775 1241.915 2008.820 ;
        RECT 1392.950 2008.760 1393.270 2008.820 ;
      LAYER via ;
        RECT 19.880 2008.760 20.140 2009.020 ;
        RECT 1392.980 2008.760 1393.240 2009.020 ;
      LAYER met2 ;
        RECT 19.880 2008.730 20.140 2009.050 ;
        RECT 1392.980 2008.730 1393.240 2009.050 ;
        RECT 19.940 1615.525 20.080 2008.730 ;
        RECT 1393.040 2000.000 1393.180 2008.730 ;
        RECT 1392.880 1999.540 1393.180 2000.000 ;
        RECT 1392.880 1996.000 1393.160 1999.540 ;
        RECT 19.870 1615.155 20.150 1615.525 ;
      LAYER via2 ;
        RECT 19.870 1615.200 20.150 1615.480 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 19.845 1615.490 20.175 1615.505 ;
        RECT -4.800 1615.190 20.175 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 19.845 1615.175 20.175 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.930 2008.620 19.250 2008.680 ;
        RECT 1400.770 2008.620 1401.090 2008.680 ;
        RECT 18.930 2008.480 1401.090 2008.620 ;
        RECT 18.930 2008.420 19.250 2008.480 ;
        RECT 1400.770 2008.420 1401.090 2008.480 ;
      LAYER via ;
        RECT 18.960 2008.420 19.220 2008.680 ;
        RECT 1400.800 2008.420 1401.060 2008.680 ;
      LAYER met2 ;
        RECT 18.960 2008.390 19.220 2008.710 ;
        RECT 1400.800 2008.390 1401.060 2008.710 ;
        RECT 19.020 1400.645 19.160 2008.390 ;
        RECT 1400.860 2000.000 1401.000 2008.390 ;
        RECT 1400.700 1999.540 1401.000 2000.000 ;
        RECT 1400.700 1996.000 1400.980 1999.540 ;
        RECT 18.950 1400.275 19.230 1400.645 ;
      LAYER via2 ;
        RECT 18.950 1400.320 19.230 1400.600 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 18.925 1400.610 19.255 1400.625 ;
        RECT -4.800 1400.310 19.255 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 18.925 1400.295 19.255 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1240.765 2008.125 1241.855 2008.295 ;
      LAYER mcon ;
        RECT 1241.685 2008.125 1241.855 2008.295 ;
      LAYER met1 ;
        RECT 18.010 2008.280 18.330 2008.340 ;
        RECT 1240.705 2008.280 1240.995 2008.325 ;
        RECT 18.010 2008.140 1240.995 2008.280 ;
        RECT 18.010 2008.080 18.330 2008.140 ;
        RECT 1240.705 2008.095 1240.995 2008.140 ;
        RECT 1241.625 2008.280 1241.915 2008.325 ;
        RECT 1408.590 2008.280 1408.910 2008.340 ;
        RECT 1241.625 2008.140 1408.910 2008.280 ;
        RECT 1241.625 2008.095 1241.915 2008.140 ;
        RECT 1408.590 2008.080 1408.910 2008.140 ;
      LAYER via ;
        RECT 18.040 2008.080 18.300 2008.340 ;
        RECT 1408.620 2008.080 1408.880 2008.340 ;
      LAYER met2 ;
        RECT 18.040 2008.050 18.300 2008.370 ;
        RECT 1408.620 2008.050 1408.880 2008.370 ;
        RECT 18.100 1185.085 18.240 2008.050 ;
        RECT 1408.680 2000.000 1408.820 2008.050 ;
        RECT 1408.520 1999.540 1408.820 2000.000 ;
        RECT 1408.520 1996.000 1408.800 1999.540 ;
        RECT 18.030 1184.715 18.310 1185.085 ;
      LAYER via2 ;
        RECT 18.030 1184.760 18.310 1185.040 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 18.005 1185.050 18.335 1185.065 ;
        RECT -4.800 1184.750 18.335 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 18.005 1184.735 18.335 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1415.050 1996.890 1415.330 1997.005 ;
        RECT 1416.340 1996.890 1416.620 2000.000 ;
        RECT 1415.050 1996.750 1416.620 1996.890 ;
        RECT 1415.050 1996.635 1415.330 1996.750 ;
        RECT 1416.340 1996.000 1416.620 1996.750 ;
        RECT 16.650 972.555 16.930 972.925 ;
        RECT 16.720 969.525 16.860 972.555 ;
        RECT 16.650 969.155 16.930 969.525 ;
      LAYER via2 ;
        RECT 1415.050 1996.680 1415.330 1996.960 ;
        RECT 16.650 972.600 16.930 972.880 ;
        RECT 16.650 969.200 16.930 969.480 ;
      LAYER met3 ;
        RECT 1414.310 1996.970 1414.690 1996.980 ;
        RECT 1415.025 1996.970 1415.355 1996.985 ;
        RECT 1414.310 1996.670 1415.355 1996.970 ;
        RECT 1414.310 1996.660 1414.690 1996.670 ;
        RECT 1415.025 1996.655 1415.355 1996.670 ;
        RECT 16.625 972.890 16.955 972.905 ;
        RECT 1414.310 972.890 1414.690 972.900 ;
        RECT 16.625 972.590 1414.690 972.890 ;
        RECT 16.625 972.575 16.955 972.590 ;
        RECT 1414.310 972.580 1414.690 972.590 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 16.625 969.490 16.955 969.505 ;
        RECT -4.800 969.190 16.955 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 16.625 969.175 16.955 969.190 ;
      LAYER via3 ;
        RECT 1414.340 1996.660 1414.660 1996.980 ;
        RECT 1414.340 972.580 1414.660 972.900 ;
      LAYER met4 ;
        RECT 1414.335 1996.655 1414.665 1996.985 ;
        RECT 1414.350 972.905 1414.650 1996.655 ;
        RECT 1414.335 972.575 1414.665 972.905 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1135.350 2005.220 1135.670 2005.280 ;
        RECT 1424.230 2005.220 1424.550 2005.280 ;
        RECT 1135.350 2005.080 1424.550 2005.220 ;
        RECT 1135.350 2005.020 1135.670 2005.080 ;
        RECT 1424.230 2005.020 1424.550 2005.080 ;
        RECT 15.710 758.780 16.030 758.840 ;
        RECT 1135.350 758.780 1135.670 758.840 ;
        RECT 15.710 758.640 1135.670 758.780 ;
        RECT 15.710 758.580 16.030 758.640 ;
        RECT 1135.350 758.580 1135.670 758.640 ;
      LAYER via ;
        RECT 1135.380 2005.020 1135.640 2005.280 ;
        RECT 1424.260 2005.020 1424.520 2005.280 ;
        RECT 15.740 758.580 16.000 758.840 ;
        RECT 1135.380 758.580 1135.640 758.840 ;
      LAYER met2 ;
        RECT 1135.380 2004.990 1135.640 2005.310 ;
        RECT 1424.260 2004.990 1424.520 2005.310 ;
        RECT 1135.440 758.870 1135.580 2004.990 ;
        RECT 1424.320 2000.000 1424.460 2004.990 ;
        RECT 1424.160 1999.540 1424.460 2000.000 ;
        RECT 1424.160 1996.000 1424.440 1999.540 ;
        RECT 15.740 758.550 16.000 758.870 ;
        RECT 1135.380 758.550 1135.640 758.870 ;
        RECT 15.800 753.965 15.940 758.550 ;
        RECT 15.730 753.595 16.010 753.965 ;
      LAYER via2 ;
        RECT 15.730 753.640 16.010 753.920 ;
      LAYER met3 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 15.705 753.930 16.035 753.945 ;
        RECT -4.800 753.630 16.035 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 15.705 753.615 16.035 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1430.690 1996.890 1430.970 1997.005 ;
        RECT 1431.980 1996.890 1432.260 2000.000 ;
        RECT 1430.690 1996.750 1432.260 1996.890 ;
        RECT 1430.690 1996.635 1430.970 1996.750 ;
        RECT 1431.980 1996.000 1432.260 1996.750 ;
        RECT 17.110 544.835 17.390 545.205 ;
        RECT 17.180 538.405 17.320 544.835 ;
        RECT 17.110 538.035 17.390 538.405 ;
      LAYER via2 ;
        RECT 1430.690 1996.680 1430.970 1996.960 ;
        RECT 17.110 544.880 17.390 545.160 ;
        RECT 17.110 538.080 17.390 538.360 ;
      LAYER met3 ;
        RECT 1428.110 1996.970 1428.490 1996.980 ;
        RECT 1430.665 1996.970 1430.995 1996.985 ;
        RECT 1428.110 1996.670 1430.995 1996.970 ;
        RECT 1428.110 1996.660 1428.490 1996.670 ;
        RECT 1430.665 1996.655 1430.995 1996.670 ;
        RECT 17.085 545.170 17.415 545.185 ;
        RECT 1428.110 545.170 1428.490 545.180 ;
        RECT 17.085 544.870 1428.490 545.170 ;
        RECT 17.085 544.855 17.415 544.870 ;
        RECT 1428.110 544.860 1428.490 544.870 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 17.085 538.370 17.415 538.385 ;
        RECT -4.800 538.070 17.415 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 17.085 538.055 17.415 538.070 ;
      LAYER via3 ;
        RECT 1428.140 1996.660 1428.460 1996.980 ;
        RECT 1428.140 544.860 1428.460 545.180 ;
      LAYER met4 ;
        RECT 1428.135 1996.655 1428.465 1996.985 ;
        RECT 1428.150 545.185 1428.450 1996.655 ;
        RECT 1428.135 544.855 1428.465 545.185 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 989.990 324.260 990.310 324.320 ;
        RECT 16.630 324.120 990.310 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 989.990 324.060 990.310 324.120 ;
      LAYER via ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 990.020 324.060 990.280 324.320 ;
      LAYER met2 ;
        RECT 1439.430 1996.890 1439.710 1997.005 ;
        RECT 1440.260 1996.890 1440.540 2000.000 ;
        RECT 1439.430 1996.750 1440.540 1996.890 ;
        RECT 1439.430 1996.635 1439.710 1996.750 ;
        RECT 1440.260 1996.000 1440.540 1996.750 ;
        RECT 990.010 1990.515 990.290 1990.885 ;
        RECT 990.080 324.350 990.220 1990.515 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 990.020 324.030 990.280 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 1439.430 1996.680 1439.710 1996.960 ;
        RECT 990.010 1990.560 990.290 1990.840 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 1439.405 1996.980 1439.735 1996.985 ;
        RECT 1439.150 1996.970 1439.735 1996.980 ;
        RECT 1438.950 1996.670 1439.735 1996.970 ;
        RECT 1439.150 1996.660 1439.735 1996.670 ;
        RECT 1439.405 1996.655 1439.735 1996.660 ;
        RECT 989.985 1990.850 990.315 1990.865 ;
        RECT 1439.150 1990.850 1439.530 1990.860 ;
        RECT 989.985 1990.550 1439.530 1990.850 ;
        RECT 989.985 1990.535 990.315 1990.550 ;
        RECT 1439.150 1990.540 1439.530 1990.550 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
      LAYER via3 ;
        RECT 1439.180 1996.660 1439.500 1996.980 ;
        RECT 1439.180 1990.540 1439.500 1990.860 ;
      LAYER met4 ;
        RECT 1439.175 1996.655 1439.505 1996.985 ;
        RECT 1439.190 1990.865 1439.490 1996.655 ;
        RECT 1439.175 1990.535 1439.505 1990.865 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1127.990 1997.740 1128.310 1997.800 ;
        RECT 1446.310 1997.740 1446.630 1997.800 ;
        RECT 1127.990 1997.600 1446.630 1997.740 ;
        RECT 1127.990 1997.540 1128.310 1997.600 ;
        RECT 1446.310 1997.540 1446.630 1997.600 ;
        RECT 15.710 110.400 16.030 110.460 ;
        RECT 1127.990 110.400 1128.310 110.460 ;
        RECT 15.710 110.260 1128.310 110.400 ;
        RECT 15.710 110.200 16.030 110.260 ;
        RECT 1127.990 110.200 1128.310 110.260 ;
      LAYER via ;
        RECT 1128.020 1997.540 1128.280 1997.800 ;
        RECT 1446.340 1997.540 1446.600 1997.800 ;
        RECT 15.740 110.200 16.000 110.460 ;
        RECT 1128.020 110.200 1128.280 110.460 ;
      LAYER met2 ;
        RECT 1128.020 1997.510 1128.280 1997.830 ;
        RECT 1446.340 1997.570 1446.600 1997.830 ;
        RECT 1448.080 1997.570 1448.360 2000.000 ;
        RECT 1446.340 1997.510 1448.360 1997.570 ;
        RECT 1128.080 110.490 1128.220 1997.510 ;
        RECT 1446.400 1997.430 1448.360 1997.510 ;
        RECT 1448.080 1996.000 1448.360 1997.430 ;
        RECT 15.740 110.170 16.000 110.490 ;
        RECT 1128.020 110.170 1128.280 110.490 ;
        RECT 15.800 107.285 15.940 110.170 ;
        RECT 15.730 106.915 16.010 107.285 ;
      LAYER via2 ;
        RECT 15.730 106.960 16.010 107.240 ;
      LAYER met3 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 15.705 107.250 16.035 107.265 ;
        RECT -4.800 106.950 16.035 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 15.705 106.935 16.035 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2466.590 2009.980 2466.910 2010.040 ;
        RECT 1179.600 2009.840 2466.910 2009.980 ;
        RECT 1179.600 2009.700 1179.740 2009.840 ;
        RECT 2466.590 2009.780 2466.910 2009.840 ;
        RECT 1179.510 2009.440 1179.830 2009.700 ;
        RECT 2466.590 855.340 2466.910 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 2466.590 855.200 2901.150 855.340 ;
        RECT 2466.590 855.140 2466.910 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 2466.620 2009.780 2466.880 2010.040 ;
        RECT 1179.540 2009.440 1179.800 2009.700 ;
        RECT 2466.620 855.140 2466.880 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 2466.620 2009.750 2466.880 2010.070 ;
        RECT 1179.540 2009.410 1179.800 2009.730 ;
        RECT 1179.600 2000.000 1179.740 2009.410 ;
        RECT 1179.440 1999.540 1179.740 2000.000 ;
        RECT 1179.440 1996.000 1179.720 1999.540 ;
        RECT 2466.680 855.430 2466.820 2009.750 ;
        RECT 2466.620 855.110 2466.880 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1187.790 2001.480 1188.110 2001.540 ;
        RECT 2066.390 2001.480 2066.710 2001.540 ;
        RECT 1187.790 2001.340 2066.710 2001.480 ;
        RECT 1187.790 2001.280 1188.110 2001.340 ;
        RECT 2066.390 2001.280 2066.710 2001.340 ;
        RECT 2066.390 1089.940 2066.710 1090.000 ;
        RECT 2900.830 1089.940 2901.150 1090.000 ;
        RECT 2066.390 1089.800 2901.150 1089.940 ;
        RECT 2066.390 1089.740 2066.710 1089.800 ;
        RECT 2900.830 1089.740 2901.150 1089.800 ;
      LAYER via ;
        RECT 1187.820 2001.280 1188.080 2001.540 ;
        RECT 2066.420 2001.280 2066.680 2001.540 ;
        RECT 2066.420 1089.740 2066.680 1090.000 ;
        RECT 2900.860 1089.740 2901.120 1090.000 ;
      LAYER met2 ;
        RECT 1187.820 2001.250 1188.080 2001.570 ;
        RECT 2066.420 2001.250 2066.680 2001.570 ;
        RECT 1187.880 2000.000 1188.020 2001.250 ;
        RECT 1187.720 1999.540 1188.020 2000.000 ;
        RECT 1187.720 1996.000 1188.000 1999.540 ;
        RECT 2066.480 1090.030 2066.620 2001.250 ;
        RECT 2066.420 1089.710 2066.680 1090.030 ;
        RECT 2900.860 1089.710 2901.120 1090.030 ;
        RECT 2900.920 1085.125 2901.060 1089.710 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
        RECT 2900.825 1085.090 2901.155 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2900.825 1084.790 2924.800 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1224.205 2009.315 1224.375 2009.655 ;
        RECT 1224.205 2009.145 1227.595 2009.315 ;
      LAYER mcon ;
        RECT 1224.205 2009.485 1224.375 2009.655 ;
        RECT 1227.425 2009.145 1227.595 2009.315 ;
      LAYER met1 ;
        RECT 1195.610 2009.640 1195.930 2009.700 ;
        RECT 1224.145 2009.640 1224.435 2009.685 ;
        RECT 1195.610 2009.500 1224.435 2009.640 ;
        RECT 1195.610 2009.440 1195.930 2009.500 ;
        RECT 1224.145 2009.455 1224.435 2009.500 ;
        RECT 1228.360 2009.500 1234.940 2009.640 ;
        RECT 1227.365 2009.300 1227.655 2009.345 ;
        RECT 1228.360 2009.300 1228.500 2009.500 ;
        RECT 1227.365 2009.160 1228.500 2009.300 ;
        RECT 1234.800 2009.300 1234.940 2009.500 ;
        RECT 2494.190 2009.300 2494.510 2009.360 ;
        RECT 1234.800 2009.160 2494.510 2009.300 ;
        RECT 1227.365 2009.115 1227.655 2009.160 ;
        RECT 2494.190 2009.100 2494.510 2009.160 ;
        RECT 2494.190 1324.540 2494.510 1324.600 ;
        RECT 2900.830 1324.540 2901.150 1324.600 ;
        RECT 2494.190 1324.400 2901.150 1324.540 ;
        RECT 2494.190 1324.340 2494.510 1324.400 ;
        RECT 2900.830 1324.340 2901.150 1324.400 ;
      LAYER via ;
        RECT 1195.640 2009.440 1195.900 2009.700 ;
        RECT 2494.220 2009.100 2494.480 2009.360 ;
        RECT 2494.220 1324.340 2494.480 1324.600 ;
        RECT 2900.860 1324.340 2901.120 1324.600 ;
      LAYER met2 ;
        RECT 1195.640 2009.410 1195.900 2009.730 ;
        RECT 1195.700 2000.000 1195.840 2009.410 ;
        RECT 2494.220 2009.070 2494.480 2009.390 ;
        RECT 1195.540 1999.540 1195.840 2000.000 ;
        RECT 1195.540 1996.000 1195.820 1999.540 ;
        RECT 2494.280 1324.630 2494.420 2009.070 ;
        RECT 2494.220 1324.310 2494.480 1324.630 ;
        RECT 2900.860 1324.310 2901.120 1324.630 ;
        RECT 2900.920 1319.725 2901.060 1324.310 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
      LAYER via2 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
      LAYER met3 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1241.685 2009.485 1241.855 2010.675 ;
      LAYER mcon ;
        RECT 1241.685 2010.505 1241.855 2010.675 ;
      LAYER met1 ;
        RECT 1203.430 2010.660 1203.750 2010.720 ;
        RECT 1241.625 2010.660 1241.915 2010.705 ;
        RECT 1203.430 2010.520 1241.915 2010.660 ;
        RECT 1203.430 2010.460 1203.750 2010.520 ;
        RECT 1241.625 2010.475 1241.915 2010.520 ;
        RECT 1241.625 2009.640 1241.915 2009.685 ;
        RECT 2501.090 2009.640 2501.410 2009.700 ;
        RECT 1241.625 2009.500 2501.410 2009.640 ;
        RECT 1241.625 2009.455 1241.915 2009.500 ;
        RECT 2501.090 2009.440 2501.410 2009.500 ;
        RECT 2501.090 1559.140 2501.410 1559.200 ;
        RECT 2900.830 1559.140 2901.150 1559.200 ;
        RECT 2501.090 1559.000 2901.150 1559.140 ;
        RECT 2501.090 1558.940 2501.410 1559.000 ;
        RECT 2900.830 1558.940 2901.150 1559.000 ;
      LAYER via ;
        RECT 1203.460 2010.460 1203.720 2010.720 ;
        RECT 2501.120 2009.440 2501.380 2009.700 ;
        RECT 2501.120 1558.940 2501.380 1559.200 ;
        RECT 2900.860 1558.940 2901.120 1559.200 ;
      LAYER met2 ;
        RECT 1203.460 2010.430 1203.720 2010.750 ;
        RECT 1203.520 2000.000 1203.660 2010.430 ;
        RECT 2501.120 2009.410 2501.380 2009.730 ;
        RECT 1203.360 1999.540 1203.660 2000.000 ;
        RECT 1203.360 1996.000 1203.640 1999.540 ;
        RECT 2501.180 1559.230 2501.320 2009.410 ;
        RECT 2501.120 1558.910 2501.380 1559.230 ;
        RECT 2900.860 1558.910 2901.120 1559.230 ;
        RECT 2900.920 1554.325 2901.060 1558.910 ;
        RECT 2900.850 1553.955 2901.130 1554.325 ;
      LAYER via2 ;
        RECT 2900.850 1554.000 2901.130 1554.280 ;
      LAYER met3 ;
        RECT 2900.825 1554.290 2901.155 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.825 1553.990 2924.800 1554.290 ;
        RECT 2900.825 1553.975 2901.155 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1631.690 1793.740 1632.010 1793.800 ;
        RECT 2900.370 1793.740 2900.690 1793.800 ;
        RECT 1631.690 1793.600 2900.690 1793.740 ;
        RECT 1631.690 1793.540 1632.010 1793.600 ;
        RECT 2900.370 1793.540 2900.690 1793.600 ;
      LAYER via ;
        RECT 1631.720 1793.540 1631.980 1793.800 ;
        RECT 2900.400 1793.540 2900.660 1793.800 ;
      LAYER met2 ;
        RECT 1211.180 1996.890 1211.460 2000.000 ;
        RECT 1212.650 1996.890 1212.930 1997.005 ;
        RECT 1211.180 1996.750 1212.930 1996.890 ;
        RECT 1211.180 1996.000 1211.460 1996.750 ;
        RECT 1212.650 1996.635 1212.930 1996.750 ;
        RECT 1631.710 1991.875 1631.990 1992.245 ;
        RECT 1631.780 1793.830 1631.920 1991.875 ;
        RECT 1631.720 1793.510 1631.980 1793.830 ;
        RECT 2900.400 1793.510 2900.660 1793.830 ;
        RECT 2900.460 1789.605 2900.600 1793.510 ;
        RECT 2900.390 1789.235 2900.670 1789.605 ;
      LAYER via2 ;
        RECT 1212.650 1996.680 1212.930 1996.960 ;
        RECT 1631.710 1991.920 1631.990 1992.200 ;
        RECT 2900.390 1789.280 2900.670 1789.560 ;
      LAYER met3 ;
        RECT 1212.625 1996.970 1212.955 1996.985 ;
        RECT 1213.750 1996.970 1214.130 1996.980 ;
        RECT 1212.625 1996.670 1214.130 1996.970 ;
        RECT 1212.625 1996.655 1212.955 1996.670 ;
        RECT 1213.750 1996.660 1214.130 1996.670 ;
        RECT 1213.750 1992.210 1214.130 1992.220 ;
        RECT 1631.685 1992.210 1632.015 1992.225 ;
        RECT 1213.750 1991.910 1632.015 1992.210 ;
        RECT 1213.750 1991.900 1214.130 1991.910 ;
        RECT 1631.685 1991.895 1632.015 1991.910 ;
        RECT 2900.365 1789.570 2900.695 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2900.365 1789.270 2924.800 1789.570 ;
        RECT 2900.365 1789.255 2900.695 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
      LAYER via3 ;
        RECT 1213.780 1996.660 1214.100 1996.980 ;
        RECT 1213.780 1991.900 1214.100 1992.220 ;
      LAYER met4 ;
        RECT 1213.775 1996.655 1214.105 1996.985 ;
        RECT 1213.790 1992.225 1214.090 1996.655 ;
        RECT 1213.775 1991.895 1214.105 1992.225 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1219.070 2021.880 1219.390 2021.940 ;
        RECT 2900.830 2021.880 2901.150 2021.940 ;
        RECT 1219.070 2021.740 2901.150 2021.880 ;
        RECT 1219.070 2021.680 1219.390 2021.740 ;
        RECT 2900.830 2021.680 2901.150 2021.740 ;
      LAYER via ;
        RECT 1219.100 2021.680 1219.360 2021.940 ;
        RECT 2900.860 2021.680 2901.120 2021.940 ;
      LAYER met2 ;
        RECT 2900.850 2023.835 2901.130 2024.205 ;
        RECT 2900.920 2021.970 2901.060 2023.835 ;
        RECT 1219.100 2021.650 1219.360 2021.970 ;
        RECT 2900.860 2021.650 2901.120 2021.970 ;
        RECT 1219.160 2000.000 1219.300 2021.650 ;
        RECT 1219.000 1999.540 1219.300 2000.000 ;
        RECT 1219.000 1996.000 1219.280 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2023.880 2901.130 2024.160 ;
      LAYER met3 ;
        RECT 2900.825 2024.170 2901.155 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2900.825 2023.870 2924.800 2024.170 ;
        RECT 2900.825 2023.855 2901.155 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1497.000 2256.680 1499.440 2256.820 ;
        RECT 1227.350 2256.480 1227.670 2256.540 ;
        RECT 1497.000 2256.480 1497.140 2256.680 ;
        RECT 1227.350 2256.340 1497.140 2256.480 ;
        RECT 1499.300 2256.480 1499.440 2256.680 ;
        RECT 2900.830 2256.480 2901.150 2256.540 ;
        RECT 1499.300 2256.340 2901.150 2256.480 ;
        RECT 1227.350 2256.280 1227.670 2256.340 ;
        RECT 2900.830 2256.280 2901.150 2256.340 ;
      LAYER via ;
        RECT 1227.380 2256.280 1227.640 2256.540 ;
        RECT 2900.860 2256.280 2901.120 2256.540 ;
      LAYER met2 ;
        RECT 2900.850 2258.435 2901.130 2258.805 ;
        RECT 2900.920 2256.570 2901.060 2258.435 ;
        RECT 1227.380 2256.250 1227.640 2256.570 ;
        RECT 2900.860 2256.250 2901.120 2256.570 ;
        RECT 1226.820 1999.610 1227.100 2000.000 ;
        RECT 1227.440 1999.610 1227.580 2256.250 ;
        RECT 1226.820 1999.470 1227.580 1999.610 ;
        RECT 1226.820 1996.000 1227.100 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 2258.480 2901.130 2258.760 ;
      LAYER met3 ;
        RECT 2900.825 2258.770 2901.155 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2900.825 2258.470 2924.800 2258.770 ;
        RECT 2900.825 2258.455 2901.155 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1179.125 1680.705 1179.295 1682.915 ;
      LAYER mcon ;
        RECT 1179.125 1682.745 1179.295 1682.915 ;
      LAYER met1 ;
        RECT 1201.590 1687.660 1201.910 1687.720 ;
        RECT 1214.930 1687.660 1215.250 1687.720 ;
        RECT 1201.590 1687.520 1215.250 1687.660 ;
        RECT 1201.590 1687.460 1201.910 1687.520 ;
        RECT 1214.930 1687.460 1215.250 1687.520 ;
        RECT 1179.065 1682.900 1179.355 1682.945 ;
        RECT 1201.590 1682.900 1201.910 1682.960 ;
        RECT 1179.065 1682.760 1201.910 1682.900 ;
        RECT 1179.065 1682.715 1179.355 1682.760 ;
        RECT 1201.590 1682.700 1201.910 1682.760 ;
        RECT 634.410 1680.860 634.730 1680.920 ;
        RECT 1179.065 1680.860 1179.355 1680.905 ;
        RECT 634.410 1680.720 1179.355 1680.860 ;
        RECT 634.410 1680.660 634.730 1680.720 ;
        RECT 1179.065 1680.675 1179.355 1680.720 ;
      LAYER via ;
        RECT 1201.620 1687.460 1201.880 1687.720 ;
        RECT 1214.960 1687.460 1215.220 1687.720 ;
        RECT 1201.620 1682.700 1201.880 1682.960 ;
        RECT 634.440 1680.660 634.700 1680.920 ;
      LAYER met2 ;
        RECT 1214.860 1700.340 1215.140 1704.000 ;
        RECT 1214.860 1700.000 1215.160 1700.340 ;
        RECT 1215.020 1687.750 1215.160 1700.000 ;
        RECT 1201.620 1687.430 1201.880 1687.750 ;
        RECT 1214.960 1687.430 1215.220 1687.750 ;
        RECT 1201.680 1682.990 1201.820 1687.430 ;
        RECT 1201.620 1682.670 1201.880 1682.990 ;
        RECT 634.440 1680.630 634.700 1680.950 ;
        RECT 634.500 17.410 634.640 1680.630 ;
        RECT 633.120 17.270 634.640 17.410 ;
        RECT 633.120 2.400 633.260 17.270 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1410.980 1690.920 1415.260 1691.060 ;
        RECT 1398.470 1690.380 1398.790 1690.440 ;
        RECT 1410.980 1690.380 1411.120 1690.920 ;
        RECT 1398.470 1690.240 1411.120 1690.380 ;
        RECT 1415.120 1690.380 1415.260 1690.920 ;
        RECT 1455.970 1690.380 1456.290 1690.440 ;
        RECT 1415.120 1690.240 1456.290 1690.380 ;
        RECT 1398.470 1690.180 1398.790 1690.240 ;
        RECT 1455.970 1690.180 1456.290 1690.240 ;
        RECT 1455.970 1680.860 1456.290 1680.920 ;
        RECT 2415.070 1680.860 2415.390 1680.920 ;
        RECT 1455.970 1680.720 2415.390 1680.860 ;
        RECT 1455.970 1680.660 1456.290 1680.720 ;
        RECT 2415.070 1680.660 2415.390 1680.720 ;
      LAYER via ;
        RECT 1398.500 1690.180 1398.760 1690.440 ;
        RECT 1456.000 1690.180 1456.260 1690.440 ;
        RECT 1456.000 1680.660 1456.260 1680.920 ;
        RECT 2415.100 1680.660 2415.360 1680.920 ;
      LAYER met2 ;
        RECT 1398.400 1700.340 1398.680 1704.000 ;
        RECT 1398.400 1700.000 1398.700 1700.340 ;
        RECT 1398.560 1690.470 1398.700 1700.000 ;
        RECT 1398.500 1690.150 1398.760 1690.470 ;
        RECT 1456.000 1690.150 1456.260 1690.470 ;
        RECT 1456.060 1680.950 1456.200 1690.150 ;
        RECT 1456.000 1680.630 1456.260 1680.950 ;
        RECT 2415.100 1680.630 2415.360 1680.950 ;
        RECT 2415.160 17.410 2415.300 1680.630 ;
        RECT 2415.160 17.270 2417.600 17.410 ;
        RECT 2417.460 2.400 2417.600 17.270 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1449.145 1687.505 1450.235 1687.675 ;
      LAYER mcon ;
        RECT 1450.065 1687.505 1450.235 1687.675 ;
      LAYER met1 ;
        RECT 1400.310 1689.020 1400.630 1689.080 ;
        RECT 1400.310 1688.880 1413.880 1689.020 ;
        RECT 1400.310 1688.820 1400.630 1688.880 ;
        RECT 1413.740 1688.000 1413.880 1688.880 ;
        RECT 1413.740 1687.860 1421.700 1688.000 ;
        RECT 1421.560 1687.660 1421.700 1687.860 ;
        RECT 1449.085 1687.660 1449.375 1687.705 ;
        RECT 1421.560 1687.520 1449.375 1687.660 ;
        RECT 1449.085 1687.475 1449.375 1687.520 ;
        RECT 1450.005 1687.660 1450.295 1687.705 ;
        RECT 1576.490 1687.660 1576.810 1687.720 ;
        RECT 1450.005 1687.520 1576.810 1687.660 ;
        RECT 1450.005 1687.475 1450.295 1687.520 ;
        RECT 1576.490 1687.460 1576.810 1687.520 ;
        RECT 1576.490 24.040 1576.810 24.100 ;
        RECT 2434.850 24.040 2435.170 24.100 ;
        RECT 1576.490 23.900 2435.170 24.040 ;
        RECT 1576.490 23.840 1576.810 23.900 ;
        RECT 2434.850 23.840 2435.170 23.900 ;
      LAYER via ;
        RECT 1400.340 1688.820 1400.600 1689.080 ;
        RECT 1576.520 1687.460 1576.780 1687.720 ;
        RECT 1576.520 23.840 1576.780 24.100 ;
        RECT 2434.880 23.840 2435.140 24.100 ;
      LAYER met2 ;
        RECT 1400.240 1700.340 1400.520 1704.000 ;
        RECT 1400.240 1700.000 1400.540 1700.340 ;
        RECT 1400.400 1689.110 1400.540 1700.000 ;
        RECT 1400.340 1688.790 1400.600 1689.110 ;
        RECT 1576.520 1687.430 1576.780 1687.750 ;
        RECT 1576.580 24.130 1576.720 1687.430 ;
        RECT 1576.520 23.810 1576.780 24.130 ;
        RECT 2434.880 23.810 2435.140 24.130 ;
        RECT 2434.940 2.400 2435.080 23.810 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1414.185 1683.765 1414.355 1686.995 ;
        RECT 1437.185 1684.445 1437.355 1688.015 ;
        RECT 1449.605 1687.845 1450.695 1688.015 ;
      LAYER mcon ;
        RECT 1437.185 1687.845 1437.355 1688.015 ;
        RECT 1450.525 1687.845 1450.695 1688.015 ;
        RECT 1414.185 1686.825 1414.355 1686.995 ;
      LAYER met1 ;
        RECT 1437.125 1688.000 1437.415 1688.045 ;
        RECT 1449.545 1688.000 1449.835 1688.045 ;
        RECT 1437.125 1687.860 1449.835 1688.000 ;
        RECT 1437.125 1687.815 1437.415 1687.860 ;
        RECT 1449.545 1687.815 1449.835 1687.860 ;
        RECT 1450.465 1688.000 1450.755 1688.045 ;
        RECT 1583.390 1688.000 1583.710 1688.060 ;
        RECT 1450.465 1687.860 1583.710 1688.000 ;
        RECT 1450.465 1687.815 1450.755 1687.860 ;
        RECT 1583.390 1687.800 1583.710 1687.860 ;
        RECT 1402.150 1686.980 1402.470 1687.040 ;
        RECT 1414.125 1686.980 1414.415 1687.025 ;
        RECT 1402.150 1686.840 1414.415 1686.980 ;
        RECT 1402.150 1686.780 1402.470 1686.840 ;
        RECT 1414.125 1686.795 1414.415 1686.840 ;
        RECT 1437.125 1684.600 1437.415 1684.645 ;
        RECT 1415.120 1684.460 1437.415 1684.600 ;
        RECT 1414.125 1683.920 1414.415 1683.965 ;
        RECT 1415.120 1683.920 1415.260 1684.460 ;
        RECT 1437.125 1684.415 1437.415 1684.460 ;
        RECT 1414.125 1683.780 1415.260 1683.920 ;
        RECT 1414.125 1683.735 1414.415 1683.780 ;
        RECT 1583.390 37.980 1583.710 38.040 ;
        RECT 2452.790 37.980 2453.110 38.040 ;
        RECT 1583.390 37.840 2453.110 37.980 ;
        RECT 1583.390 37.780 1583.710 37.840 ;
        RECT 2452.790 37.780 2453.110 37.840 ;
      LAYER via ;
        RECT 1583.420 1687.800 1583.680 1688.060 ;
        RECT 1402.180 1686.780 1402.440 1687.040 ;
        RECT 1583.420 37.780 1583.680 38.040 ;
        RECT 2452.820 37.780 2453.080 38.040 ;
      LAYER met2 ;
        RECT 1402.080 1700.340 1402.360 1704.000 ;
        RECT 1402.080 1700.000 1402.380 1700.340 ;
        RECT 1402.240 1687.070 1402.380 1700.000 ;
        RECT 1583.420 1687.770 1583.680 1688.090 ;
        RECT 1402.180 1686.750 1402.440 1687.070 ;
        RECT 1583.480 38.070 1583.620 1687.770 ;
        RECT 1583.420 37.750 1583.680 38.070 ;
        RECT 2452.820 37.750 2453.080 38.070 ;
        RECT 2452.880 2.400 2453.020 37.750 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1447.765 1688.525 1448.855 1688.695 ;
        RECT 1449.145 1688.525 1451.155 1688.695 ;
        RECT 1450.985 1686.485 1451.155 1688.525 ;
        RECT 1494.225 1686.485 1494.395 1689.375 ;
      LAYER mcon ;
        RECT 1494.225 1689.205 1494.395 1689.375 ;
        RECT 1448.685 1688.525 1448.855 1688.695 ;
      LAYER met1 ;
        RECT 1494.165 1689.360 1494.455 1689.405 ;
        RECT 1514.390 1689.360 1514.710 1689.420 ;
        RECT 1494.165 1689.220 1514.710 1689.360 ;
        RECT 1494.165 1689.175 1494.455 1689.220 ;
        RECT 1514.390 1689.160 1514.710 1689.220 ;
        RECT 1447.690 1688.680 1448.010 1688.740 ;
        RECT 1448.625 1688.680 1448.915 1688.725 ;
        RECT 1449.085 1688.680 1449.375 1688.725 ;
        RECT 1447.690 1688.540 1448.205 1688.680 ;
        RECT 1448.625 1688.540 1449.375 1688.680 ;
        RECT 1447.690 1688.480 1448.010 1688.540 ;
        RECT 1448.625 1688.495 1448.915 1688.540 ;
        RECT 1449.085 1688.495 1449.375 1688.540 ;
        RECT 1450.925 1686.640 1451.215 1686.685 ;
        RECT 1494.165 1686.640 1494.455 1686.685 ;
        RECT 1450.925 1686.500 1494.455 1686.640 ;
        RECT 1450.925 1686.455 1451.215 1686.500 ;
        RECT 1494.165 1686.455 1494.455 1686.500 ;
        RECT 1514.390 44.780 1514.710 44.840 ;
        RECT 2470.730 44.780 2471.050 44.840 ;
        RECT 1514.390 44.640 2471.050 44.780 ;
        RECT 1514.390 44.580 1514.710 44.640 ;
        RECT 2470.730 44.580 2471.050 44.640 ;
      LAYER via ;
        RECT 1514.420 1689.160 1514.680 1689.420 ;
        RECT 1447.720 1688.480 1447.980 1688.740 ;
        RECT 1514.420 44.580 1514.680 44.840 ;
        RECT 2470.760 44.580 2471.020 44.840 ;
      LAYER met2 ;
        RECT 1403.920 1700.340 1404.200 1704.000 ;
        RECT 1403.920 1700.000 1404.220 1700.340 ;
        RECT 1404.080 1689.645 1404.220 1700.000 ;
        RECT 1404.010 1689.275 1404.290 1689.645 ;
        RECT 1447.710 1689.275 1447.990 1689.645 ;
        RECT 1447.780 1688.770 1447.920 1689.275 ;
        RECT 1514.420 1689.130 1514.680 1689.450 ;
        RECT 1447.720 1688.450 1447.980 1688.770 ;
        RECT 1514.480 44.870 1514.620 1689.130 ;
        RECT 1514.420 44.550 1514.680 44.870 ;
        RECT 2470.760 44.550 2471.020 44.870 ;
        RECT 2470.820 2.400 2470.960 44.550 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
      LAYER via2 ;
        RECT 1404.010 1689.320 1404.290 1689.600 ;
        RECT 1447.710 1689.320 1447.990 1689.600 ;
      LAYER met3 ;
        RECT 1403.985 1689.610 1404.315 1689.625 ;
        RECT 1447.685 1689.610 1448.015 1689.625 ;
        RECT 1403.985 1689.310 1448.015 1689.610 ;
        RECT 1403.985 1689.295 1404.315 1689.310 ;
        RECT 1447.685 1689.295 1448.015 1689.310 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1412.805 1689.885 1413.895 1690.055 ;
        RECT 1413.725 1684.785 1413.895 1689.885 ;
        RECT 1457.425 1685.125 1457.595 1686.995 ;
        RECT 1544.825 1686.825 1545.455 1686.995 ;
        RECT 1545.285 1686.485 1545.455 1686.825 ;
        RECT 1607.845 1686.655 1608.015 1686.995 ;
        RECT 1559.085 1686.485 1560.175 1686.655 ;
        RECT 1607.385 1686.485 1608.015 1686.655 ;
        RECT 1642.345 1685.805 1642.515 1686.655 ;
        RECT 1690.645 1685.125 1690.815 1685.975 ;
        RECT 1738.485 1685.125 1738.655 1686.655 ;
        RECT 1738.945 1685.805 1739.115 1686.655 ;
        RECT 1760.565 1685.805 1760.735 1686.655 ;
        RECT 1787.245 1685.805 1787.415 1686.655 ;
        RECT 1835.085 1685.805 1835.255 1686.655 ;
        RECT 1835.545 1685.805 1835.715 1686.655 ;
        RECT 1857.165 1685.805 1857.335 1686.655 ;
        RECT 1883.845 1685.805 1884.015 1686.655 ;
        RECT 1931.685 1685.805 1931.855 1686.655 ;
        RECT 1932.145 1685.805 1932.315 1686.655 ;
        RECT 1953.765 1685.805 1953.935 1686.655 ;
        RECT 1980.445 1685.805 1980.615 1686.655 ;
        RECT 2028.285 1685.805 2028.455 1686.655 ;
        RECT 2028.745 1685.805 2028.915 1686.655 ;
        RECT 2050.365 1685.805 2050.535 1686.655 ;
        RECT 2077.045 1685.805 2077.215 1686.655 ;
        RECT 2124.885 1685.805 2125.055 1686.655 ;
        RECT 2125.345 1685.805 2125.515 1686.655 ;
        RECT 2146.965 1685.805 2147.135 1686.655 ;
        RECT 2173.645 1685.805 2173.815 1686.655 ;
        RECT 2221.485 1685.805 2221.655 1686.655 ;
        RECT 2221.945 1685.805 2222.115 1686.655 ;
        RECT 2243.565 1685.805 2243.735 1686.655 ;
        RECT 2270.245 1685.805 2270.415 1686.655 ;
        RECT 2318.085 1685.805 2318.255 1686.655 ;
        RECT 2318.545 1685.805 2318.715 1686.655 ;
        RECT 2340.165 1685.805 2340.335 1686.655 ;
        RECT 2366.845 1685.805 2367.015 1686.655 ;
        RECT 2414.685 1685.805 2414.855 1686.995 ;
        RECT 2417.905 1683.425 2418.075 1686.995 ;
      LAYER mcon ;
        RECT 1457.425 1686.825 1457.595 1686.995 ;
        RECT 1607.845 1686.825 1608.015 1686.995 ;
        RECT 2414.685 1686.825 2414.855 1686.995 ;
        RECT 1560.005 1686.485 1560.175 1686.655 ;
        RECT 1642.345 1686.485 1642.515 1686.655 ;
        RECT 1738.485 1686.485 1738.655 1686.655 ;
        RECT 1690.645 1685.805 1690.815 1685.975 ;
        RECT 1738.945 1686.485 1739.115 1686.655 ;
        RECT 1760.565 1686.485 1760.735 1686.655 ;
        RECT 1787.245 1686.485 1787.415 1686.655 ;
        RECT 1835.085 1686.485 1835.255 1686.655 ;
        RECT 1835.545 1686.485 1835.715 1686.655 ;
        RECT 1857.165 1686.485 1857.335 1686.655 ;
        RECT 1883.845 1686.485 1884.015 1686.655 ;
        RECT 1931.685 1686.485 1931.855 1686.655 ;
        RECT 1932.145 1686.485 1932.315 1686.655 ;
        RECT 1953.765 1686.485 1953.935 1686.655 ;
        RECT 1980.445 1686.485 1980.615 1686.655 ;
        RECT 2028.285 1686.485 2028.455 1686.655 ;
        RECT 2028.745 1686.485 2028.915 1686.655 ;
        RECT 2050.365 1686.485 2050.535 1686.655 ;
        RECT 2077.045 1686.485 2077.215 1686.655 ;
        RECT 2124.885 1686.485 2125.055 1686.655 ;
        RECT 2125.345 1686.485 2125.515 1686.655 ;
        RECT 2146.965 1686.485 2147.135 1686.655 ;
        RECT 2173.645 1686.485 2173.815 1686.655 ;
        RECT 2221.485 1686.485 2221.655 1686.655 ;
        RECT 2221.945 1686.485 2222.115 1686.655 ;
        RECT 2243.565 1686.485 2243.735 1686.655 ;
        RECT 2270.245 1686.485 2270.415 1686.655 ;
        RECT 2318.085 1686.485 2318.255 1686.655 ;
        RECT 2318.545 1686.485 2318.715 1686.655 ;
        RECT 2340.165 1686.485 2340.335 1686.655 ;
        RECT 2366.845 1686.485 2367.015 1686.655 ;
        RECT 2417.905 1686.825 2418.075 1686.995 ;
      LAYER met1 ;
        RECT 1405.830 1690.040 1406.150 1690.100 ;
        RECT 1412.745 1690.040 1413.035 1690.085 ;
        RECT 1405.830 1689.900 1413.035 1690.040 ;
        RECT 1405.830 1689.840 1406.150 1689.900 ;
        RECT 1412.745 1689.855 1413.035 1689.900 ;
        RECT 1457.365 1686.980 1457.655 1687.025 ;
        RECT 1544.765 1686.980 1545.055 1687.025 ;
        RECT 1457.365 1686.840 1545.055 1686.980 ;
        RECT 1457.365 1686.795 1457.655 1686.840 ;
        RECT 1544.765 1686.795 1545.055 1686.840 ;
        RECT 1607.785 1686.980 1608.075 1687.025 ;
        RECT 2414.625 1686.980 2414.915 1687.025 ;
        RECT 2417.845 1686.980 2418.135 1687.025 ;
        RECT 1607.785 1686.840 1642.500 1686.980 ;
        RECT 1607.785 1686.795 1608.075 1686.840 ;
        RECT 1642.360 1686.685 1642.500 1686.840 ;
        RECT 1738.500 1686.840 1739.100 1686.980 ;
        RECT 1738.500 1686.685 1738.640 1686.840 ;
        RECT 1738.960 1686.685 1739.100 1686.840 ;
        RECT 1835.100 1686.840 1835.700 1686.980 ;
        RECT 1835.100 1686.685 1835.240 1686.840 ;
        RECT 1835.560 1686.685 1835.700 1686.840 ;
        RECT 1931.700 1686.840 1932.300 1686.980 ;
        RECT 1931.700 1686.685 1931.840 1686.840 ;
        RECT 1932.160 1686.685 1932.300 1686.840 ;
        RECT 2028.300 1686.840 2028.900 1686.980 ;
        RECT 2028.300 1686.685 2028.440 1686.840 ;
        RECT 2028.760 1686.685 2028.900 1686.840 ;
        RECT 2124.900 1686.840 2125.500 1686.980 ;
        RECT 2124.900 1686.685 2125.040 1686.840 ;
        RECT 2125.360 1686.685 2125.500 1686.840 ;
        RECT 2221.500 1686.840 2222.100 1686.980 ;
        RECT 2221.500 1686.685 2221.640 1686.840 ;
        RECT 2221.960 1686.685 2222.100 1686.840 ;
        RECT 2318.100 1686.840 2318.700 1686.980 ;
        RECT 2318.100 1686.685 2318.240 1686.840 ;
        RECT 2318.560 1686.685 2318.700 1686.840 ;
        RECT 2414.625 1686.840 2418.135 1686.980 ;
        RECT 2414.625 1686.795 2414.915 1686.840 ;
        RECT 2417.845 1686.795 2418.135 1686.840 ;
        RECT 1545.225 1686.640 1545.515 1686.685 ;
        RECT 1559.025 1686.640 1559.315 1686.685 ;
        RECT 1545.225 1686.500 1559.315 1686.640 ;
        RECT 1545.225 1686.455 1545.515 1686.500 ;
        RECT 1559.025 1686.455 1559.315 1686.500 ;
        RECT 1559.945 1686.640 1560.235 1686.685 ;
        RECT 1607.325 1686.640 1607.615 1686.685 ;
        RECT 1559.945 1686.500 1607.615 1686.640 ;
        RECT 1559.945 1686.455 1560.235 1686.500 ;
        RECT 1607.325 1686.455 1607.615 1686.500 ;
        RECT 1642.285 1686.455 1642.575 1686.685 ;
        RECT 1738.425 1686.455 1738.715 1686.685 ;
        RECT 1738.885 1686.455 1739.175 1686.685 ;
        RECT 1760.505 1686.640 1760.795 1686.685 ;
        RECT 1787.185 1686.640 1787.475 1686.685 ;
        RECT 1760.505 1686.500 1787.475 1686.640 ;
        RECT 1760.505 1686.455 1760.795 1686.500 ;
        RECT 1787.185 1686.455 1787.475 1686.500 ;
        RECT 1835.025 1686.455 1835.315 1686.685 ;
        RECT 1835.485 1686.455 1835.775 1686.685 ;
        RECT 1857.105 1686.640 1857.395 1686.685 ;
        RECT 1883.785 1686.640 1884.075 1686.685 ;
        RECT 1857.105 1686.500 1884.075 1686.640 ;
        RECT 1857.105 1686.455 1857.395 1686.500 ;
        RECT 1883.785 1686.455 1884.075 1686.500 ;
        RECT 1931.625 1686.455 1931.915 1686.685 ;
        RECT 1932.085 1686.455 1932.375 1686.685 ;
        RECT 1953.705 1686.640 1953.995 1686.685 ;
        RECT 1980.385 1686.640 1980.675 1686.685 ;
        RECT 1953.705 1686.500 1980.675 1686.640 ;
        RECT 1953.705 1686.455 1953.995 1686.500 ;
        RECT 1980.385 1686.455 1980.675 1686.500 ;
        RECT 2028.225 1686.455 2028.515 1686.685 ;
        RECT 2028.685 1686.455 2028.975 1686.685 ;
        RECT 2050.305 1686.640 2050.595 1686.685 ;
        RECT 2076.985 1686.640 2077.275 1686.685 ;
        RECT 2050.305 1686.500 2077.275 1686.640 ;
        RECT 2050.305 1686.455 2050.595 1686.500 ;
        RECT 2076.985 1686.455 2077.275 1686.500 ;
        RECT 2124.825 1686.455 2125.115 1686.685 ;
        RECT 2125.285 1686.455 2125.575 1686.685 ;
        RECT 2146.905 1686.640 2147.195 1686.685 ;
        RECT 2173.585 1686.640 2173.875 1686.685 ;
        RECT 2146.905 1686.500 2173.875 1686.640 ;
        RECT 2146.905 1686.455 2147.195 1686.500 ;
        RECT 2173.585 1686.455 2173.875 1686.500 ;
        RECT 2221.425 1686.455 2221.715 1686.685 ;
        RECT 2221.885 1686.455 2222.175 1686.685 ;
        RECT 2243.505 1686.640 2243.795 1686.685 ;
        RECT 2270.185 1686.640 2270.475 1686.685 ;
        RECT 2243.505 1686.500 2270.475 1686.640 ;
        RECT 2243.505 1686.455 2243.795 1686.500 ;
        RECT 2270.185 1686.455 2270.475 1686.500 ;
        RECT 2318.025 1686.455 2318.315 1686.685 ;
        RECT 2318.485 1686.455 2318.775 1686.685 ;
        RECT 2340.105 1686.640 2340.395 1686.685 ;
        RECT 2366.785 1686.640 2367.075 1686.685 ;
        RECT 2340.105 1686.500 2367.075 1686.640 ;
        RECT 2340.105 1686.455 2340.395 1686.500 ;
        RECT 2366.785 1686.455 2367.075 1686.500 ;
        RECT 1642.285 1685.960 1642.575 1686.005 ;
        RECT 1690.585 1685.960 1690.875 1686.005 ;
        RECT 1642.285 1685.820 1690.875 1685.960 ;
        RECT 1642.285 1685.775 1642.575 1685.820 ;
        RECT 1690.585 1685.775 1690.875 1685.820 ;
        RECT 1738.885 1685.960 1739.175 1686.005 ;
        RECT 1760.505 1685.960 1760.795 1686.005 ;
        RECT 1738.885 1685.820 1760.795 1685.960 ;
        RECT 1738.885 1685.775 1739.175 1685.820 ;
        RECT 1760.505 1685.775 1760.795 1685.820 ;
        RECT 1787.185 1685.960 1787.475 1686.005 ;
        RECT 1835.025 1685.960 1835.315 1686.005 ;
        RECT 1787.185 1685.820 1835.315 1685.960 ;
        RECT 1787.185 1685.775 1787.475 1685.820 ;
        RECT 1835.025 1685.775 1835.315 1685.820 ;
        RECT 1835.485 1685.960 1835.775 1686.005 ;
        RECT 1857.105 1685.960 1857.395 1686.005 ;
        RECT 1835.485 1685.820 1857.395 1685.960 ;
        RECT 1835.485 1685.775 1835.775 1685.820 ;
        RECT 1857.105 1685.775 1857.395 1685.820 ;
        RECT 1883.785 1685.960 1884.075 1686.005 ;
        RECT 1931.625 1685.960 1931.915 1686.005 ;
        RECT 1883.785 1685.820 1931.915 1685.960 ;
        RECT 1883.785 1685.775 1884.075 1685.820 ;
        RECT 1931.625 1685.775 1931.915 1685.820 ;
        RECT 1932.085 1685.960 1932.375 1686.005 ;
        RECT 1953.705 1685.960 1953.995 1686.005 ;
        RECT 1932.085 1685.820 1953.995 1685.960 ;
        RECT 1932.085 1685.775 1932.375 1685.820 ;
        RECT 1953.705 1685.775 1953.995 1685.820 ;
        RECT 1980.385 1685.960 1980.675 1686.005 ;
        RECT 2028.225 1685.960 2028.515 1686.005 ;
        RECT 1980.385 1685.820 2028.515 1685.960 ;
        RECT 1980.385 1685.775 1980.675 1685.820 ;
        RECT 2028.225 1685.775 2028.515 1685.820 ;
        RECT 2028.685 1685.960 2028.975 1686.005 ;
        RECT 2050.305 1685.960 2050.595 1686.005 ;
        RECT 2028.685 1685.820 2050.595 1685.960 ;
        RECT 2028.685 1685.775 2028.975 1685.820 ;
        RECT 2050.305 1685.775 2050.595 1685.820 ;
        RECT 2076.985 1685.960 2077.275 1686.005 ;
        RECT 2124.825 1685.960 2125.115 1686.005 ;
        RECT 2076.985 1685.820 2125.115 1685.960 ;
        RECT 2076.985 1685.775 2077.275 1685.820 ;
        RECT 2124.825 1685.775 2125.115 1685.820 ;
        RECT 2125.285 1685.960 2125.575 1686.005 ;
        RECT 2146.905 1685.960 2147.195 1686.005 ;
        RECT 2125.285 1685.820 2147.195 1685.960 ;
        RECT 2125.285 1685.775 2125.575 1685.820 ;
        RECT 2146.905 1685.775 2147.195 1685.820 ;
        RECT 2173.585 1685.960 2173.875 1686.005 ;
        RECT 2221.425 1685.960 2221.715 1686.005 ;
        RECT 2173.585 1685.820 2221.715 1685.960 ;
        RECT 2173.585 1685.775 2173.875 1685.820 ;
        RECT 2221.425 1685.775 2221.715 1685.820 ;
        RECT 2221.885 1685.960 2222.175 1686.005 ;
        RECT 2243.505 1685.960 2243.795 1686.005 ;
        RECT 2221.885 1685.820 2243.795 1685.960 ;
        RECT 2221.885 1685.775 2222.175 1685.820 ;
        RECT 2243.505 1685.775 2243.795 1685.820 ;
        RECT 2270.185 1685.960 2270.475 1686.005 ;
        RECT 2318.025 1685.960 2318.315 1686.005 ;
        RECT 2270.185 1685.820 2318.315 1685.960 ;
        RECT 2270.185 1685.775 2270.475 1685.820 ;
        RECT 2318.025 1685.775 2318.315 1685.820 ;
        RECT 2318.485 1685.960 2318.775 1686.005 ;
        RECT 2340.105 1685.960 2340.395 1686.005 ;
        RECT 2318.485 1685.820 2340.395 1685.960 ;
        RECT 2318.485 1685.775 2318.775 1685.820 ;
        RECT 2340.105 1685.775 2340.395 1685.820 ;
        RECT 2366.785 1685.960 2367.075 1686.005 ;
        RECT 2414.625 1685.960 2414.915 1686.005 ;
        RECT 2366.785 1685.820 2414.915 1685.960 ;
        RECT 2366.785 1685.775 2367.075 1685.820 ;
        RECT 2414.625 1685.775 2414.915 1685.820 ;
        RECT 1457.365 1685.280 1457.655 1685.325 ;
        RECT 1438.580 1685.140 1457.655 1685.280 ;
        RECT 1413.665 1684.940 1413.955 1684.985 ;
        RECT 1438.580 1684.940 1438.720 1685.140 ;
        RECT 1457.365 1685.095 1457.655 1685.140 ;
        RECT 1690.585 1685.280 1690.875 1685.325 ;
        RECT 1738.425 1685.280 1738.715 1685.325 ;
        RECT 1690.585 1685.140 1738.715 1685.280 ;
        RECT 1690.585 1685.095 1690.875 1685.140 ;
        RECT 1738.425 1685.095 1738.715 1685.140 ;
        RECT 1413.665 1684.800 1438.720 1684.940 ;
        RECT 1413.665 1684.755 1413.955 1684.800 ;
        RECT 2417.845 1683.580 2418.135 1683.625 ;
        RECT 2445.890 1683.580 2446.210 1683.640 ;
        RECT 2417.845 1683.440 2446.210 1683.580 ;
        RECT 2417.845 1683.395 2418.135 1683.440 ;
        RECT 2445.890 1683.380 2446.210 1683.440 ;
        RECT 2445.890 24.040 2446.210 24.100 ;
        RECT 2488.670 24.040 2488.990 24.100 ;
        RECT 2445.890 23.900 2488.990 24.040 ;
        RECT 2445.890 23.840 2446.210 23.900 ;
        RECT 2488.670 23.840 2488.990 23.900 ;
      LAYER via ;
        RECT 1405.860 1689.840 1406.120 1690.100 ;
        RECT 2445.920 1683.380 2446.180 1683.640 ;
        RECT 2445.920 23.840 2446.180 24.100 ;
        RECT 2488.700 23.840 2488.960 24.100 ;
      LAYER met2 ;
        RECT 1405.760 1700.340 1406.040 1704.000 ;
        RECT 1405.760 1700.000 1406.060 1700.340 ;
        RECT 1405.920 1690.130 1406.060 1700.000 ;
        RECT 1405.860 1689.810 1406.120 1690.130 ;
        RECT 2445.920 1683.350 2446.180 1683.670 ;
        RECT 2445.980 24.130 2446.120 1683.350 ;
        RECT 2445.920 23.810 2446.180 24.130 ;
        RECT 2488.700 23.810 2488.960 24.130 ;
        RECT 2488.760 2.400 2488.900 23.810 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1422.925 1685.465 1423.095 1686.655 ;
        RECT 1450.525 1673.565 1450.695 1686.655 ;
      LAYER mcon ;
        RECT 1422.925 1686.485 1423.095 1686.655 ;
        RECT 1450.525 1686.485 1450.695 1686.655 ;
      LAYER met1 ;
        RECT 1422.865 1686.640 1423.155 1686.685 ;
        RECT 1450.465 1686.640 1450.755 1686.685 ;
        RECT 1422.865 1686.500 1450.755 1686.640 ;
        RECT 1422.865 1686.455 1423.155 1686.500 ;
        RECT 1450.465 1686.455 1450.755 1686.500 ;
        RECT 1407.670 1685.960 1407.990 1686.020 ;
        RECT 1407.670 1685.820 1412.960 1685.960 ;
        RECT 1407.670 1685.760 1407.990 1685.820 ;
        RECT 1412.820 1685.620 1412.960 1685.820 ;
        RECT 1422.865 1685.620 1423.155 1685.665 ;
        RECT 1412.820 1685.480 1423.155 1685.620 ;
        RECT 1422.865 1685.435 1423.155 1685.480 ;
        RECT 1450.465 1673.720 1450.755 1673.765 ;
        RECT 2504.770 1673.720 2505.090 1673.780 ;
        RECT 1450.465 1673.580 2505.090 1673.720 ;
        RECT 1450.465 1673.535 1450.755 1673.580 ;
        RECT 2504.770 1673.520 2505.090 1673.580 ;
      LAYER via ;
        RECT 1407.700 1685.760 1407.960 1686.020 ;
        RECT 2504.800 1673.520 2505.060 1673.780 ;
      LAYER met2 ;
        RECT 1407.600 1700.340 1407.880 1704.000 ;
        RECT 1407.600 1700.000 1407.900 1700.340 ;
        RECT 1407.760 1686.050 1407.900 1700.000 ;
        RECT 1407.700 1685.730 1407.960 1686.050 ;
        RECT 2504.800 1673.490 2505.060 1673.810 ;
        RECT 2504.860 17.410 2505.000 1673.490 ;
        RECT 2504.860 17.270 2506.380 17.410 ;
        RECT 2506.240 2.400 2506.380 17.270 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1449.605 1688.865 1450.235 1689.035 ;
      LAYER mcon ;
        RECT 1450.065 1688.865 1450.235 1689.035 ;
      LAYER met1 ;
        RECT 1438.490 1689.020 1438.810 1689.080 ;
        RECT 1449.545 1689.020 1449.835 1689.065 ;
        RECT 1438.490 1688.880 1449.835 1689.020 ;
        RECT 1438.490 1688.820 1438.810 1688.880 ;
        RECT 1449.545 1688.835 1449.835 1688.880 ;
        RECT 1450.005 1689.020 1450.295 1689.065 ;
        RECT 1507.490 1689.020 1507.810 1689.080 ;
        RECT 1450.005 1688.880 1507.810 1689.020 ;
        RECT 1450.005 1688.835 1450.295 1688.880 ;
        RECT 1507.490 1688.820 1507.810 1688.880 ;
        RECT 1507.490 58.720 1507.810 58.780 ;
        RECT 2518.570 58.720 2518.890 58.780 ;
        RECT 1507.490 58.580 2518.890 58.720 ;
        RECT 1507.490 58.520 1507.810 58.580 ;
        RECT 2518.570 58.520 2518.890 58.580 ;
      LAYER via ;
        RECT 1438.520 1688.820 1438.780 1689.080 ;
        RECT 1507.520 1688.820 1507.780 1689.080 ;
        RECT 1507.520 58.520 1507.780 58.780 ;
        RECT 2518.600 58.520 2518.860 58.780 ;
      LAYER met2 ;
        RECT 1409.440 1700.340 1409.720 1704.000 ;
        RECT 1409.440 1700.000 1409.740 1700.340 ;
        RECT 1409.600 1688.965 1409.740 1700.000 ;
        RECT 1438.520 1688.965 1438.780 1689.110 ;
        RECT 1409.530 1688.595 1409.810 1688.965 ;
        RECT 1438.510 1688.595 1438.790 1688.965 ;
        RECT 1507.520 1688.790 1507.780 1689.110 ;
        RECT 1507.580 58.810 1507.720 1688.790 ;
        RECT 1507.520 58.490 1507.780 58.810 ;
        RECT 2518.600 58.490 2518.860 58.810 ;
        RECT 2518.660 17.410 2518.800 58.490 ;
        RECT 2518.660 17.270 2524.320 17.410 ;
        RECT 2524.180 2.400 2524.320 17.270 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
      LAYER via2 ;
        RECT 1409.530 1688.640 1409.810 1688.920 ;
        RECT 1438.510 1688.640 1438.790 1688.920 ;
      LAYER met3 ;
        RECT 1409.505 1688.930 1409.835 1688.945 ;
        RECT 1438.485 1688.930 1438.815 1688.945 ;
        RECT 1409.505 1688.630 1438.815 1688.930 ;
        RECT 1409.505 1688.615 1409.835 1688.630 ;
        RECT 1438.485 1688.615 1438.815 1688.630 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1414.645 1690.225 1415.275 1690.395 ;
        RECT 1415.105 1688.865 1415.275 1690.225 ;
        RECT 1437.645 1685.975 1437.815 1689.035 ;
        RECT 1437.645 1685.805 1439.655 1685.975 ;
      LAYER mcon ;
        RECT 1437.645 1688.865 1437.815 1689.035 ;
        RECT 1439.485 1685.805 1439.655 1685.975 ;
      LAYER met1 ;
        RECT 1411.350 1690.380 1411.670 1690.440 ;
        RECT 1414.585 1690.380 1414.875 1690.425 ;
        RECT 1411.350 1690.240 1414.875 1690.380 ;
        RECT 1411.350 1690.180 1411.670 1690.240 ;
        RECT 1414.585 1690.195 1414.875 1690.240 ;
        RECT 1415.045 1689.020 1415.335 1689.065 ;
        RECT 1437.585 1689.020 1437.875 1689.065 ;
        RECT 1415.045 1688.880 1437.875 1689.020 ;
        RECT 1415.045 1688.835 1415.335 1688.880 ;
        RECT 1437.585 1688.835 1437.875 1688.880 ;
        RECT 1439.425 1685.960 1439.715 1686.005 ;
        RECT 1459.190 1685.960 1459.510 1686.020 ;
        RECT 1439.425 1685.820 1459.510 1685.960 ;
        RECT 1439.425 1685.775 1439.715 1685.820 ;
        RECT 1459.190 1685.760 1459.510 1685.820 ;
        RECT 1459.190 65.520 1459.510 65.580 ;
        RECT 2539.270 65.520 2539.590 65.580 ;
        RECT 1459.190 65.380 2539.590 65.520 ;
        RECT 1459.190 65.320 1459.510 65.380 ;
        RECT 2539.270 65.320 2539.590 65.380 ;
      LAYER via ;
        RECT 1411.380 1690.180 1411.640 1690.440 ;
        RECT 1459.220 1685.760 1459.480 1686.020 ;
        RECT 1459.220 65.320 1459.480 65.580 ;
        RECT 2539.300 65.320 2539.560 65.580 ;
      LAYER met2 ;
        RECT 1411.280 1700.340 1411.560 1704.000 ;
        RECT 1411.280 1700.000 1411.580 1700.340 ;
        RECT 1411.440 1690.470 1411.580 1700.000 ;
        RECT 1411.380 1690.150 1411.640 1690.470 ;
        RECT 1459.220 1685.730 1459.480 1686.050 ;
        RECT 1459.280 65.610 1459.420 1685.730 ;
        RECT 1459.220 65.290 1459.480 65.610 ;
        RECT 2539.300 65.290 2539.560 65.610 ;
        RECT 2539.360 17.410 2539.500 65.290 ;
        RECT 2539.360 17.270 2542.260 17.410 ;
        RECT 2542.120 2.400 2542.260 17.270 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1440.330 1689.360 1440.650 1689.420 ;
        RECT 1493.690 1689.360 1494.010 1689.420 ;
        RECT 1440.330 1689.220 1494.010 1689.360 ;
        RECT 1440.330 1689.160 1440.650 1689.220 ;
        RECT 1493.690 1689.160 1494.010 1689.220 ;
        RECT 1493.690 72.320 1494.010 72.380 ;
        RECT 2560.430 72.320 2560.750 72.380 ;
        RECT 1493.690 72.180 2560.750 72.320 ;
        RECT 1493.690 72.120 1494.010 72.180 ;
        RECT 2560.430 72.120 2560.750 72.180 ;
      LAYER via ;
        RECT 1440.360 1689.160 1440.620 1689.420 ;
        RECT 1493.720 1689.160 1493.980 1689.420 ;
        RECT 1493.720 72.120 1493.980 72.380 ;
        RECT 2560.460 72.120 2560.720 72.380 ;
      LAYER met2 ;
        RECT 1413.120 1700.340 1413.400 1704.000 ;
        RECT 1413.120 1700.000 1413.420 1700.340 ;
        RECT 1413.280 1690.325 1413.420 1700.000 ;
        RECT 1413.210 1689.955 1413.490 1690.325 ;
        RECT 1440.350 1689.955 1440.630 1690.325 ;
        RECT 1440.420 1689.450 1440.560 1689.955 ;
        RECT 1440.360 1689.130 1440.620 1689.450 ;
        RECT 1493.720 1689.130 1493.980 1689.450 ;
        RECT 1493.780 72.410 1493.920 1689.130 ;
        RECT 1493.720 72.090 1493.980 72.410 ;
        RECT 2560.460 72.090 2560.720 72.410 ;
        RECT 2560.520 7.210 2560.660 72.090 ;
        RECT 2560.060 7.070 2560.660 7.210 ;
        RECT 2560.060 2.400 2560.200 7.070 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
      LAYER via2 ;
        RECT 1413.210 1690.000 1413.490 1690.280 ;
        RECT 1440.350 1690.000 1440.630 1690.280 ;
      LAYER met3 ;
        RECT 1413.185 1690.290 1413.515 1690.305 ;
        RECT 1440.325 1690.290 1440.655 1690.305 ;
        RECT 1413.185 1689.990 1440.655 1690.290 ;
        RECT 1413.185 1689.975 1413.515 1689.990 ;
        RECT 1440.325 1689.975 1440.655 1689.990 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1434.885 1689.545 1435.055 1690.735 ;
        RECT 1439.945 1686.145 1440.115 1690.735 ;
      LAYER mcon ;
        RECT 1434.885 1690.565 1435.055 1690.735 ;
        RECT 1439.945 1690.565 1440.115 1690.735 ;
      LAYER met1 ;
        RECT 1434.825 1690.720 1435.115 1690.765 ;
        RECT 1439.885 1690.720 1440.175 1690.765 ;
        RECT 1434.825 1690.580 1440.175 1690.720 ;
        RECT 1434.825 1690.535 1435.115 1690.580 ;
        RECT 1439.885 1690.535 1440.175 1690.580 ;
        RECT 1415.030 1689.700 1415.350 1689.760 ;
        RECT 1434.825 1689.700 1435.115 1689.745 ;
        RECT 1415.030 1689.560 1435.115 1689.700 ;
        RECT 1415.030 1689.500 1415.350 1689.560 ;
        RECT 1434.825 1689.515 1435.115 1689.560 ;
        RECT 1439.885 1686.300 1440.175 1686.345 ;
        RECT 1452.290 1686.300 1452.610 1686.360 ;
        RECT 1439.885 1686.160 1452.610 1686.300 ;
        RECT 1439.885 1686.115 1440.175 1686.160 ;
        RECT 1452.290 1686.100 1452.610 1686.160 ;
        RECT 1452.290 79.460 1452.610 79.520 ;
        RECT 2573.770 79.460 2574.090 79.520 ;
        RECT 1452.290 79.320 2574.090 79.460 ;
        RECT 1452.290 79.260 1452.610 79.320 ;
        RECT 2573.770 79.260 2574.090 79.320 ;
      LAYER via ;
        RECT 1415.060 1689.500 1415.320 1689.760 ;
        RECT 1452.320 1686.100 1452.580 1686.360 ;
        RECT 1452.320 79.260 1452.580 79.520 ;
        RECT 2573.800 79.260 2574.060 79.520 ;
      LAYER met2 ;
        RECT 1414.960 1700.340 1415.240 1704.000 ;
        RECT 1414.960 1700.000 1415.260 1700.340 ;
        RECT 1415.120 1689.790 1415.260 1700.000 ;
        RECT 1415.060 1689.470 1415.320 1689.790 ;
        RECT 1452.320 1686.070 1452.580 1686.390 ;
        RECT 1452.380 79.550 1452.520 1686.070 ;
        RECT 1452.320 79.230 1452.580 79.550 ;
        RECT 2573.800 79.230 2574.060 79.550 ;
        RECT 2573.860 17.410 2574.000 79.230 ;
        RECT 2573.860 17.270 2578.140 17.410 ;
        RECT 2578.000 2.400 2578.140 17.270 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1201.130 1689.360 1201.450 1689.420 ;
        RECT 1232.870 1689.360 1233.190 1689.420 ;
        RECT 1201.130 1689.220 1233.190 1689.360 ;
        RECT 1201.130 1689.160 1201.450 1689.220 ;
        RECT 1232.870 1689.160 1233.190 1689.220 ;
        RECT 813.810 1674.060 814.130 1674.120 ;
        RECT 1201.130 1674.060 1201.450 1674.120 ;
        RECT 813.810 1673.920 1201.450 1674.060 ;
        RECT 813.810 1673.860 814.130 1673.920 ;
        RECT 1201.130 1673.860 1201.450 1673.920 ;
      LAYER via ;
        RECT 1201.160 1689.160 1201.420 1689.420 ;
        RECT 1232.900 1689.160 1233.160 1689.420 ;
        RECT 813.840 1673.860 814.100 1674.120 ;
        RECT 1201.160 1673.860 1201.420 1674.120 ;
      LAYER met2 ;
        RECT 1232.800 1700.340 1233.080 1704.000 ;
        RECT 1232.800 1700.000 1233.100 1700.340 ;
        RECT 1232.960 1689.450 1233.100 1700.000 ;
        RECT 1201.160 1689.130 1201.420 1689.450 ;
        RECT 1232.900 1689.130 1233.160 1689.450 ;
        RECT 1201.220 1674.150 1201.360 1689.130 ;
        RECT 813.840 1673.830 814.100 1674.150 ;
        RECT 1201.160 1673.830 1201.420 1674.150 ;
        RECT 813.900 17.410 814.040 1673.830 ;
        RECT 811.600 17.270 814.040 17.410 ;
        RECT 811.600 2.400 811.740 17.270 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1416.870 1685.960 1417.190 1686.020 ;
        RECT 1420.090 1685.960 1420.410 1686.020 ;
        RECT 1416.870 1685.820 1420.410 1685.960 ;
        RECT 1416.870 1685.760 1417.190 1685.820 ;
        RECT 1420.090 1685.760 1420.410 1685.820 ;
        RECT 1420.090 1678.280 1420.410 1678.540 ;
        RECT 1420.180 1677.800 1420.320 1678.280 ;
        RECT 1420.180 1677.660 1421.240 1677.800 ;
        RECT 1421.100 1677.520 1421.240 1677.660 ;
        RECT 1421.010 1677.260 1421.330 1677.520 ;
        RECT 1421.010 1666.580 1421.330 1666.640 ;
        RECT 2594.470 1666.580 2594.790 1666.640 ;
        RECT 1421.010 1666.440 2594.790 1666.580 ;
        RECT 1421.010 1666.380 1421.330 1666.440 ;
        RECT 2594.470 1666.380 2594.790 1666.440 ;
      LAYER via ;
        RECT 1416.900 1685.760 1417.160 1686.020 ;
        RECT 1420.120 1685.760 1420.380 1686.020 ;
        RECT 1420.120 1678.280 1420.380 1678.540 ;
        RECT 1421.040 1677.260 1421.300 1677.520 ;
        RECT 1421.040 1666.380 1421.300 1666.640 ;
        RECT 2594.500 1666.380 2594.760 1666.640 ;
      LAYER met2 ;
        RECT 1416.800 1700.340 1417.080 1704.000 ;
        RECT 1416.800 1700.000 1417.100 1700.340 ;
        RECT 1416.960 1686.050 1417.100 1700.000 ;
        RECT 1416.900 1685.730 1417.160 1686.050 ;
        RECT 1420.120 1685.730 1420.380 1686.050 ;
        RECT 1420.180 1678.570 1420.320 1685.730 ;
        RECT 1420.120 1678.250 1420.380 1678.570 ;
        RECT 1421.040 1677.230 1421.300 1677.550 ;
        RECT 1421.100 1666.670 1421.240 1677.230 ;
        RECT 1421.040 1666.350 1421.300 1666.670 ;
        RECT 2594.500 1666.350 2594.760 1666.670 ;
        RECT 2594.560 17.410 2594.700 1666.350 ;
        RECT 2594.560 17.270 2595.620 17.410 ;
        RECT 2595.480 2.400 2595.620 17.270 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1418.710 1687.660 1419.030 1687.720 ;
        RECT 1420.550 1687.660 1420.870 1687.720 ;
        RECT 1418.710 1687.520 1420.870 1687.660 ;
        RECT 1418.710 1687.460 1419.030 1687.520 ;
        RECT 1420.550 1687.460 1420.870 1687.520 ;
        RECT 1420.550 1680.520 1420.870 1680.580 ;
        RECT 2608.270 1680.520 2608.590 1680.580 ;
        RECT 1420.550 1680.380 2608.590 1680.520 ;
        RECT 1420.550 1680.320 1420.870 1680.380 ;
        RECT 2608.270 1680.320 2608.590 1680.380 ;
      LAYER via ;
        RECT 1418.740 1687.460 1419.000 1687.720 ;
        RECT 1420.580 1687.460 1420.840 1687.720 ;
        RECT 1420.580 1680.320 1420.840 1680.580 ;
        RECT 2608.300 1680.320 2608.560 1680.580 ;
      LAYER met2 ;
        RECT 1418.640 1700.340 1418.920 1704.000 ;
        RECT 1418.640 1700.000 1418.940 1700.340 ;
        RECT 1418.800 1687.750 1418.940 1700.000 ;
        RECT 1418.740 1687.430 1419.000 1687.750 ;
        RECT 1420.580 1687.430 1420.840 1687.750 ;
        RECT 1420.640 1680.610 1420.780 1687.430 ;
        RECT 1420.580 1680.290 1420.840 1680.610 ;
        RECT 2608.300 1680.290 2608.560 1680.610 ;
        RECT 2608.360 17.410 2608.500 1680.290 ;
        RECT 2608.360 17.270 2613.560 17.410 ;
        RECT 2613.420 2.400 2613.560 17.270 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1439.485 1689.205 1439.655 1690.055 ;
      LAYER mcon ;
        RECT 1439.485 1689.885 1439.655 1690.055 ;
      LAYER met1 ;
        RECT 1439.425 1690.040 1439.715 1690.085 ;
        RECT 1486.790 1690.040 1487.110 1690.100 ;
        RECT 1439.425 1689.900 1487.110 1690.040 ;
        RECT 1439.425 1689.855 1439.715 1689.900 ;
        RECT 1486.790 1689.840 1487.110 1689.900 ;
        RECT 1420.550 1689.360 1420.870 1689.420 ;
        RECT 1439.425 1689.360 1439.715 1689.405 ;
        RECT 1420.550 1689.220 1439.715 1689.360 ;
        RECT 1420.550 1689.160 1420.870 1689.220 ;
        RECT 1439.425 1689.175 1439.715 1689.220 ;
        RECT 1486.790 93.060 1487.110 93.120 ;
        RECT 2628.970 93.060 2629.290 93.120 ;
        RECT 1486.790 92.920 2629.290 93.060 ;
        RECT 1486.790 92.860 1487.110 92.920 ;
        RECT 2628.970 92.860 2629.290 92.920 ;
      LAYER via ;
        RECT 1486.820 1689.840 1487.080 1690.100 ;
        RECT 1420.580 1689.160 1420.840 1689.420 ;
        RECT 1486.820 92.860 1487.080 93.120 ;
        RECT 2629.000 92.860 2629.260 93.120 ;
      LAYER met2 ;
        RECT 1420.480 1700.340 1420.760 1704.000 ;
        RECT 1420.480 1700.000 1420.780 1700.340 ;
        RECT 1420.640 1689.450 1420.780 1700.000 ;
        RECT 1486.820 1689.810 1487.080 1690.130 ;
        RECT 1420.580 1689.130 1420.840 1689.450 ;
        RECT 1486.880 93.150 1487.020 1689.810 ;
        RECT 1486.820 92.830 1487.080 93.150 ;
        RECT 2629.000 92.830 2629.260 93.150 ;
        RECT 2629.060 17.410 2629.200 92.830 ;
        RECT 2629.060 17.270 2631.500 17.410 ;
        RECT 2631.360 2.400 2631.500 17.270 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1427.065 1684.105 1427.235 1688.355 ;
      LAYER mcon ;
        RECT 1427.065 1688.185 1427.235 1688.355 ;
      LAYER met1 ;
        RECT 1422.390 1688.340 1422.710 1688.400 ;
        RECT 1427.005 1688.340 1427.295 1688.385 ;
        RECT 1422.390 1688.200 1427.295 1688.340 ;
        RECT 1422.390 1688.140 1422.710 1688.200 ;
        RECT 1427.005 1688.155 1427.295 1688.200 ;
        RECT 1426.990 1684.260 1427.310 1684.320 ;
        RECT 1426.795 1684.120 1427.310 1684.260 ;
        RECT 1426.990 1684.060 1427.310 1684.120 ;
        RECT 1426.990 1659.780 1427.310 1659.840 ;
        RECT 2642.770 1659.780 2643.090 1659.840 ;
        RECT 1426.990 1659.640 2643.090 1659.780 ;
        RECT 1426.990 1659.580 1427.310 1659.640 ;
        RECT 2642.770 1659.580 2643.090 1659.640 ;
        RECT 2642.770 16.900 2643.090 16.960 ;
        RECT 2649.210 16.900 2649.530 16.960 ;
        RECT 2642.770 16.760 2649.530 16.900 ;
        RECT 2642.770 16.700 2643.090 16.760 ;
        RECT 2649.210 16.700 2649.530 16.760 ;
      LAYER via ;
        RECT 1422.420 1688.140 1422.680 1688.400 ;
        RECT 1427.020 1684.060 1427.280 1684.320 ;
        RECT 1427.020 1659.580 1427.280 1659.840 ;
        RECT 2642.800 1659.580 2643.060 1659.840 ;
        RECT 2642.800 16.700 2643.060 16.960 ;
        RECT 2649.240 16.700 2649.500 16.960 ;
      LAYER met2 ;
        RECT 1422.320 1700.340 1422.600 1704.000 ;
        RECT 1422.320 1700.000 1422.620 1700.340 ;
        RECT 1422.480 1688.430 1422.620 1700.000 ;
        RECT 1422.420 1688.110 1422.680 1688.430 ;
        RECT 1427.020 1684.030 1427.280 1684.350 ;
        RECT 1427.080 1659.870 1427.220 1684.030 ;
        RECT 1427.020 1659.550 1427.280 1659.870 ;
        RECT 2642.800 1659.550 2643.060 1659.870 ;
        RECT 2642.860 16.990 2643.000 1659.550 ;
        RECT 2642.800 16.670 2643.060 16.990 ;
        RECT 2649.240 16.670 2649.500 16.990 ;
        RECT 2649.300 2.400 2649.440 16.670 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1424.230 1688.000 1424.550 1688.060 ;
        RECT 1427.450 1688.000 1427.770 1688.060 ;
        RECT 1424.230 1687.860 1427.770 1688.000 ;
        RECT 1424.230 1687.800 1424.550 1687.860 ;
        RECT 1427.450 1687.800 1427.770 1687.860 ;
        RECT 1427.450 1673.380 1427.770 1673.440 ;
        RECT 2663.470 1673.380 2663.790 1673.440 ;
        RECT 1427.450 1673.240 2663.790 1673.380 ;
        RECT 1427.450 1673.180 1427.770 1673.240 ;
        RECT 2663.470 1673.180 2663.790 1673.240 ;
      LAYER via ;
        RECT 1424.260 1687.800 1424.520 1688.060 ;
        RECT 1427.480 1687.800 1427.740 1688.060 ;
        RECT 1427.480 1673.180 1427.740 1673.440 ;
        RECT 2663.500 1673.180 2663.760 1673.440 ;
      LAYER met2 ;
        RECT 1424.160 1700.340 1424.440 1704.000 ;
        RECT 1424.160 1700.000 1424.460 1700.340 ;
        RECT 1424.320 1688.090 1424.460 1700.000 ;
        RECT 1424.260 1687.770 1424.520 1688.090 ;
        RECT 1427.480 1687.770 1427.740 1688.090 ;
        RECT 1427.540 1673.470 1427.680 1687.770 ;
        RECT 1427.480 1673.150 1427.740 1673.470 ;
        RECT 2663.500 1673.150 2663.760 1673.470 ;
        RECT 2663.560 17.410 2663.700 1673.150 ;
        RECT 2663.560 17.270 2667.380 17.410 ;
        RECT 2667.240 2.400 2667.380 17.270 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1427.910 1652.640 1428.230 1652.700 ;
        RECT 2684.170 1652.640 2684.490 1652.700 ;
        RECT 1427.910 1652.500 2684.490 1652.640 ;
        RECT 1427.910 1652.440 1428.230 1652.500 ;
        RECT 2684.170 1652.440 2684.490 1652.500 ;
      LAYER via ;
        RECT 1427.940 1652.440 1428.200 1652.700 ;
        RECT 2684.200 1652.440 2684.460 1652.700 ;
      LAYER met2 ;
        RECT 1426.000 1700.340 1426.280 1704.000 ;
        RECT 1426.000 1700.000 1426.300 1700.340 ;
        RECT 1426.160 1684.885 1426.300 1700.000 ;
        RECT 1426.090 1684.515 1426.370 1684.885 ;
        RECT 1427.930 1684.515 1428.210 1684.885 ;
        RECT 1428.000 1652.730 1428.140 1684.515 ;
        RECT 1427.940 1652.410 1428.200 1652.730 ;
        RECT 2684.200 1652.410 2684.460 1652.730 ;
        RECT 2684.260 17.410 2684.400 1652.410 ;
        RECT 2684.260 17.270 2684.860 17.410 ;
        RECT 2684.720 2.400 2684.860 17.270 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
      LAYER via2 ;
        RECT 1426.090 1684.560 1426.370 1684.840 ;
        RECT 1427.930 1684.560 1428.210 1684.840 ;
      LAYER met3 ;
        RECT 1426.065 1684.850 1426.395 1684.865 ;
        RECT 1427.905 1684.850 1428.235 1684.865 ;
        RECT 1426.065 1684.550 1428.235 1684.850 ;
        RECT 1426.065 1684.535 1426.395 1684.550 ;
        RECT 1427.905 1684.535 1428.235 1684.550 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1427.985 1645.345 1428.155 1685.295 ;
      LAYER mcon ;
        RECT 1427.985 1685.125 1428.155 1685.295 ;
      LAYER met1 ;
        RECT 1427.910 1685.280 1428.230 1685.340 ;
        RECT 1427.715 1685.140 1428.230 1685.280 ;
        RECT 1427.910 1685.080 1428.230 1685.140 ;
        RECT 1427.925 1645.500 1428.215 1645.545 ;
        RECT 2697.970 1645.500 2698.290 1645.560 ;
        RECT 1427.925 1645.360 2698.290 1645.500 ;
        RECT 1427.925 1645.315 1428.215 1645.360 ;
        RECT 2697.970 1645.300 2698.290 1645.360 ;
      LAYER via ;
        RECT 1427.940 1685.080 1428.200 1685.340 ;
        RECT 2698.000 1645.300 2698.260 1645.560 ;
      LAYER met2 ;
        RECT 1427.840 1700.340 1428.120 1704.000 ;
        RECT 1427.840 1700.000 1428.140 1700.340 ;
        RECT 1428.000 1685.370 1428.140 1700.000 ;
        RECT 1427.940 1685.050 1428.200 1685.370 ;
        RECT 2698.000 1645.270 2698.260 1645.590 ;
        RECT 2698.060 17.410 2698.200 1645.270 ;
        RECT 2698.060 17.270 2702.800 17.410 ;
        RECT 2702.660 2.400 2702.800 17.270 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1449.145 1683.425 1449.315 1686.995 ;
      LAYER mcon ;
        RECT 1449.145 1686.825 1449.315 1686.995 ;
      LAYER met1 ;
        RECT 1429.750 1686.980 1430.070 1687.040 ;
        RECT 1449.085 1686.980 1449.375 1687.025 ;
        RECT 1429.750 1686.840 1449.375 1686.980 ;
        RECT 1429.750 1686.780 1430.070 1686.840 ;
        RECT 1449.085 1686.795 1449.375 1686.840 ;
        RECT 1449.085 1683.580 1449.375 1683.625 ;
        RECT 1473.450 1683.580 1473.770 1683.640 ;
        RECT 1449.085 1683.440 1473.770 1683.580 ;
        RECT 1449.085 1683.395 1449.375 1683.440 ;
        RECT 1473.450 1683.380 1473.770 1683.440 ;
        RECT 1473.450 99.860 1473.770 99.920 ;
        RECT 2718.670 99.860 2718.990 99.920 ;
        RECT 1473.450 99.720 2718.990 99.860 ;
        RECT 1473.450 99.660 1473.770 99.720 ;
        RECT 2718.670 99.660 2718.990 99.720 ;
      LAYER via ;
        RECT 1429.780 1686.780 1430.040 1687.040 ;
        RECT 1473.480 1683.380 1473.740 1683.640 ;
        RECT 1473.480 99.660 1473.740 99.920 ;
        RECT 2718.700 99.660 2718.960 99.920 ;
      LAYER met2 ;
        RECT 1429.680 1700.340 1429.960 1704.000 ;
        RECT 1429.680 1700.000 1429.980 1700.340 ;
        RECT 1429.840 1687.070 1429.980 1700.000 ;
        RECT 1429.780 1686.750 1430.040 1687.070 ;
        RECT 1473.480 1683.350 1473.740 1683.670 ;
        RECT 1473.540 99.950 1473.680 1683.350 ;
        RECT 1473.480 99.630 1473.740 99.950 ;
        RECT 2718.700 99.630 2718.960 99.950 ;
        RECT 2718.760 17.410 2718.900 99.630 ;
        RECT 2718.760 17.270 2720.740 17.410 ;
        RECT 2720.600 2.400 2720.740 17.270 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1431.590 1685.280 1431.910 1685.340 ;
        RECT 1434.810 1685.280 1435.130 1685.340 ;
        RECT 1431.590 1685.140 1435.130 1685.280 ;
        RECT 1431.590 1685.080 1431.910 1685.140 ;
        RECT 1434.810 1685.080 1435.130 1685.140 ;
        RECT 1434.810 1666.240 1435.130 1666.300 ;
        RECT 2732.470 1666.240 2732.790 1666.300 ;
        RECT 1434.810 1666.100 2732.790 1666.240 ;
        RECT 1434.810 1666.040 1435.130 1666.100 ;
        RECT 2732.470 1666.040 2732.790 1666.100 ;
        RECT 2732.470 18.260 2732.790 18.320 ;
        RECT 2738.450 18.260 2738.770 18.320 ;
        RECT 2732.470 18.120 2738.770 18.260 ;
        RECT 2732.470 18.060 2732.790 18.120 ;
        RECT 2738.450 18.060 2738.770 18.120 ;
      LAYER via ;
        RECT 1431.620 1685.080 1431.880 1685.340 ;
        RECT 1434.840 1685.080 1435.100 1685.340 ;
        RECT 1434.840 1666.040 1435.100 1666.300 ;
        RECT 2732.500 1666.040 2732.760 1666.300 ;
        RECT 2732.500 18.060 2732.760 18.320 ;
        RECT 2738.480 18.060 2738.740 18.320 ;
      LAYER met2 ;
        RECT 1431.520 1700.340 1431.800 1704.000 ;
        RECT 1431.520 1700.000 1431.820 1700.340 ;
        RECT 1431.680 1685.370 1431.820 1700.000 ;
        RECT 1431.620 1685.050 1431.880 1685.370 ;
        RECT 1434.840 1685.050 1435.100 1685.370 ;
        RECT 1434.900 1666.330 1435.040 1685.050 ;
        RECT 1434.840 1666.010 1435.100 1666.330 ;
        RECT 2732.500 1666.010 2732.760 1666.330 ;
        RECT 2732.560 18.350 2732.700 1666.010 ;
        RECT 2732.500 18.030 2732.760 18.350 ;
        RECT 2738.480 18.030 2738.740 18.350 ;
        RECT 2738.540 2.400 2738.680 18.030 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1433.430 1638.700 1433.750 1638.760 ;
        RECT 2753.170 1638.700 2753.490 1638.760 ;
        RECT 1433.430 1638.560 2753.490 1638.700 ;
        RECT 1433.430 1638.500 1433.750 1638.560 ;
        RECT 2753.170 1638.500 2753.490 1638.560 ;
      LAYER via ;
        RECT 1433.460 1638.500 1433.720 1638.760 ;
        RECT 2753.200 1638.500 2753.460 1638.760 ;
      LAYER met2 ;
        RECT 1433.360 1700.340 1433.640 1704.000 ;
        RECT 1433.360 1700.000 1433.660 1700.340 ;
        RECT 1433.520 1638.790 1433.660 1700.000 ;
        RECT 1433.460 1638.470 1433.720 1638.790 ;
        RECT 2753.200 1638.470 2753.460 1638.790 ;
        RECT 2753.260 17.410 2753.400 1638.470 ;
        RECT 2753.260 17.270 2756.160 17.410 ;
        RECT 2756.020 2.400 2756.160 17.270 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1179.585 1686.485 1179.755 1688.015 ;
      LAYER mcon ;
        RECT 1179.585 1687.845 1179.755 1688.015 ;
      LAYER met1 ;
        RECT 1179.525 1688.000 1179.815 1688.045 ;
        RECT 1234.710 1688.000 1235.030 1688.060 ;
        RECT 1179.525 1687.860 1235.030 1688.000 ;
        RECT 1179.525 1687.815 1179.815 1687.860 ;
        RECT 1234.710 1687.800 1235.030 1687.860 ;
        RECT 1134.890 1686.640 1135.210 1686.700 ;
        RECT 1179.525 1686.640 1179.815 1686.685 ;
        RECT 1134.890 1686.500 1179.815 1686.640 ;
        RECT 1134.890 1686.440 1135.210 1686.500 ;
        RECT 1179.525 1686.455 1179.815 1686.500 ;
        RECT 834.510 58.720 834.830 58.780 ;
        RECT 1134.890 58.720 1135.210 58.780 ;
        RECT 834.510 58.580 1135.210 58.720 ;
        RECT 834.510 58.520 834.830 58.580 ;
        RECT 1134.890 58.520 1135.210 58.580 ;
      LAYER via ;
        RECT 1234.740 1687.800 1235.000 1688.060 ;
        RECT 1134.920 1686.440 1135.180 1686.700 ;
        RECT 834.540 58.520 834.800 58.780 ;
        RECT 1134.920 58.520 1135.180 58.780 ;
      LAYER met2 ;
        RECT 1234.640 1700.340 1234.920 1704.000 ;
        RECT 1234.640 1700.000 1234.940 1700.340 ;
        RECT 1234.800 1688.090 1234.940 1700.000 ;
        RECT 1234.740 1687.770 1235.000 1688.090 ;
        RECT 1134.920 1686.410 1135.180 1686.730 ;
        RECT 1134.980 58.810 1135.120 1686.410 ;
        RECT 834.540 58.490 834.800 58.810 ;
        RECT 1134.920 58.490 1135.180 58.810 ;
        RECT 834.600 17.410 834.740 58.490 ;
        RECT 829.540 17.270 834.740 17.410 ;
        RECT 829.540 2.400 829.680 17.270 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1449.145 1689.545 1450.695 1689.715 ;
      LAYER mcon ;
        RECT 1450.525 1689.545 1450.695 1689.715 ;
      LAYER met1 ;
        RECT 1435.270 1690.040 1435.590 1690.100 ;
        RECT 1435.270 1689.900 1439.180 1690.040 ;
        RECT 1435.270 1689.840 1435.590 1689.900 ;
        RECT 1439.040 1689.700 1439.180 1689.900 ;
        RECT 1449.085 1689.700 1449.375 1689.745 ;
        RECT 1439.040 1689.560 1449.375 1689.700 ;
        RECT 1449.085 1689.515 1449.375 1689.560 ;
        RECT 1450.465 1689.700 1450.755 1689.745 ;
        RECT 1454.130 1689.700 1454.450 1689.760 ;
        RECT 1450.465 1689.560 1454.450 1689.700 ;
        RECT 1450.465 1689.515 1450.755 1689.560 ;
        RECT 1454.130 1689.500 1454.450 1689.560 ;
        RECT 1454.130 1631.900 1454.450 1631.960 ;
        RECT 2773.870 1631.900 2774.190 1631.960 ;
        RECT 1454.130 1631.760 2774.190 1631.900 ;
        RECT 1454.130 1631.700 1454.450 1631.760 ;
        RECT 2773.870 1631.700 2774.190 1631.760 ;
      LAYER via ;
        RECT 1435.300 1689.840 1435.560 1690.100 ;
        RECT 1454.160 1689.500 1454.420 1689.760 ;
        RECT 1454.160 1631.700 1454.420 1631.960 ;
        RECT 2773.900 1631.700 2774.160 1631.960 ;
      LAYER met2 ;
        RECT 1435.200 1700.340 1435.480 1704.000 ;
        RECT 1435.200 1700.000 1435.500 1700.340 ;
        RECT 1435.360 1690.130 1435.500 1700.000 ;
        RECT 1435.300 1689.810 1435.560 1690.130 ;
        RECT 1454.160 1689.470 1454.420 1689.790 ;
        RECT 1454.220 1631.990 1454.360 1689.470 ;
        RECT 1454.160 1631.670 1454.420 1631.990 ;
        RECT 2773.900 1631.670 2774.160 1631.990 ;
        RECT 2773.960 2.400 2774.100 1631.670 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1437.110 1685.960 1437.430 1686.020 ;
        RECT 1438.950 1685.960 1439.270 1686.020 ;
        RECT 1437.110 1685.820 1439.270 1685.960 ;
        RECT 1437.110 1685.760 1437.430 1685.820 ;
        RECT 1438.950 1685.760 1439.270 1685.820 ;
        RECT 1438.950 1680.180 1439.270 1680.240 ;
        RECT 2787.670 1680.180 2787.990 1680.240 ;
        RECT 1438.950 1680.040 2787.990 1680.180 ;
        RECT 1438.950 1679.980 1439.270 1680.040 ;
        RECT 2787.670 1679.980 2787.990 1680.040 ;
      LAYER via ;
        RECT 1437.140 1685.760 1437.400 1686.020 ;
        RECT 1438.980 1685.760 1439.240 1686.020 ;
        RECT 1438.980 1679.980 1439.240 1680.240 ;
        RECT 2787.700 1679.980 2787.960 1680.240 ;
      LAYER met2 ;
        RECT 1437.040 1700.340 1437.320 1704.000 ;
        RECT 1437.040 1700.000 1437.340 1700.340 ;
        RECT 1437.200 1686.050 1437.340 1700.000 ;
        RECT 1437.140 1685.730 1437.400 1686.050 ;
        RECT 1438.980 1685.730 1439.240 1686.050 ;
        RECT 1439.040 1680.270 1439.180 1685.730 ;
        RECT 1438.980 1679.950 1439.240 1680.270 ;
        RECT 2787.700 1679.950 2787.960 1680.270 ;
        RECT 2787.760 17.410 2787.900 1679.950 ;
        RECT 2787.760 17.270 2792.040 17.410 ;
        RECT 2791.900 2.400 2792.040 17.270 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1438.950 1688.340 1439.270 1688.400 ;
        RECT 1604.090 1688.340 1604.410 1688.400 ;
        RECT 1438.950 1688.200 1604.410 1688.340 ;
        RECT 1438.950 1688.140 1439.270 1688.200 ;
        RECT 1604.090 1688.140 1604.410 1688.200 ;
        RECT 1604.090 107.000 1604.410 107.060 ;
        RECT 2808.370 107.000 2808.690 107.060 ;
        RECT 1604.090 106.860 2808.690 107.000 ;
        RECT 1604.090 106.800 1604.410 106.860 ;
        RECT 2808.370 106.800 2808.690 106.860 ;
      LAYER via ;
        RECT 1438.980 1688.140 1439.240 1688.400 ;
        RECT 1604.120 1688.140 1604.380 1688.400 ;
        RECT 1604.120 106.800 1604.380 107.060 ;
        RECT 2808.400 106.800 2808.660 107.060 ;
      LAYER met2 ;
        RECT 1438.880 1700.340 1439.160 1704.000 ;
        RECT 1438.880 1700.000 1439.180 1700.340 ;
        RECT 1439.040 1688.430 1439.180 1700.000 ;
        RECT 1438.980 1688.110 1439.240 1688.430 ;
        RECT 1604.120 1688.110 1604.380 1688.430 ;
        RECT 1604.180 107.090 1604.320 1688.110 ;
        RECT 1604.120 106.770 1604.380 107.090 ;
        RECT 2808.400 106.770 2808.660 107.090 ;
        RECT 2808.460 17.410 2808.600 106.770 ;
        RECT 2808.460 17.270 2809.980 17.410 ;
        RECT 2809.840 2.400 2809.980 17.270 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1440.790 1624.760 1441.110 1624.820 ;
        RECT 2822.170 1624.760 2822.490 1624.820 ;
        RECT 1440.790 1624.620 2822.490 1624.760 ;
        RECT 1440.790 1624.560 1441.110 1624.620 ;
        RECT 2822.170 1624.560 2822.490 1624.620 ;
      LAYER via ;
        RECT 1440.820 1624.560 1441.080 1624.820 ;
        RECT 2822.200 1624.560 2822.460 1624.820 ;
      LAYER met2 ;
        RECT 1440.720 1700.340 1441.000 1704.000 ;
        RECT 1440.720 1700.000 1441.020 1700.340 ;
        RECT 1440.880 1624.850 1441.020 1700.000 ;
        RECT 1440.820 1624.530 1441.080 1624.850 ;
        RECT 2822.200 1624.530 2822.460 1624.850 ;
        RECT 2822.260 17.410 2822.400 1624.530 ;
        RECT 2822.260 17.270 2827.920 17.410 ;
        RECT 2827.780 2.400 2827.920 17.270 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1442.630 1684.940 1442.950 1685.000 ;
        RECT 1453.670 1684.940 1453.990 1685.000 ;
        RECT 1442.630 1684.800 1453.990 1684.940 ;
        RECT 1442.630 1684.740 1442.950 1684.800 ;
        RECT 1453.670 1684.740 1453.990 1684.800 ;
        RECT 1453.670 1617.960 1453.990 1618.020 ;
        RECT 2842.870 1617.960 2843.190 1618.020 ;
        RECT 1453.670 1617.820 2843.190 1617.960 ;
        RECT 1453.670 1617.760 1453.990 1617.820 ;
        RECT 2842.870 1617.760 2843.190 1617.820 ;
      LAYER via ;
        RECT 1442.660 1684.740 1442.920 1685.000 ;
        RECT 1453.700 1684.740 1453.960 1685.000 ;
        RECT 1453.700 1617.760 1453.960 1618.020 ;
        RECT 2842.900 1617.760 2843.160 1618.020 ;
      LAYER met2 ;
        RECT 1442.560 1700.340 1442.840 1704.000 ;
        RECT 1442.560 1700.000 1442.860 1700.340 ;
        RECT 1442.720 1685.030 1442.860 1700.000 ;
        RECT 1442.660 1684.710 1442.920 1685.030 ;
        RECT 1453.700 1684.710 1453.960 1685.030 ;
        RECT 1453.760 1618.050 1453.900 1684.710 ;
        RECT 1453.700 1617.730 1453.960 1618.050 ;
        RECT 2842.900 1617.730 2843.160 1618.050 ;
        RECT 2842.960 16.730 2843.100 1617.730 ;
        RECT 2842.960 16.590 2845.400 16.730 ;
        RECT 2845.260 2.400 2845.400 16.590 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1444.470 1684.260 1444.790 1684.320 ;
        RECT 1453.210 1684.260 1453.530 1684.320 ;
        RECT 1444.470 1684.120 1453.530 1684.260 ;
        RECT 1444.470 1684.060 1444.790 1684.120 ;
        RECT 1453.210 1684.060 1453.530 1684.120 ;
        RECT 1453.210 1604.360 1453.530 1604.420 ;
        RECT 2857.130 1604.360 2857.450 1604.420 ;
        RECT 1453.210 1604.220 2857.450 1604.360 ;
        RECT 1453.210 1604.160 1453.530 1604.220 ;
        RECT 2857.130 1604.160 2857.450 1604.220 ;
        RECT 2857.130 18.600 2857.450 18.660 ;
        RECT 2863.110 18.600 2863.430 18.660 ;
        RECT 2857.130 18.460 2863.430 18.600 ;
        RECT 2857.130 18.400 2857.450 18.460 ;
        RECT 2863.110 18.400 2863.430 18.460 ;
      LAYER via ;
        RECT 1444.500 1684.060 1444.760 1684.320 ;
        RECT 1453.240 1684.060 1453.500 1684.320 ;
        RECT 1453.240 1604.160 1453.500 1604.420 ;
        RECT 2857.160 1604.160 2857.420 1604.420 ;
        RECT 2857.160 18.400 2857.420 18.660 ;
        RECT 2863.140 18.400 2863.400 18.660 ;
      LAYER met2 ;
        RECT 1444.400 1700.340 1444.680 1704.000 ;
        RECT 1444.400 1700.000 1444.700 1700.340 ;
        RECT 1444.560 1684.350 1444.700 1700.000 ;
        RECT 1444.500 1684.030 1444.760 1684.350 ;
        RECT 1453.240 1684.030 1453.500 1684.350 ;
        RECT 1453.300 1604.450 1453.440 1684.030 ;
        RECT 1453.240 1604.130 1453.500 1604.450 ;
        RECT 2857.160 1604.130 2857.420 1604.450 ;
        RECT 2857.220 18.690 2857.360 1604.130 ;
        RECT 2857.160 18.370 2857.420 18.690 ;
        RECT 2863.140 18.370 2863.400 18.690 ;
        RECT 2863.200 2.400 2863.340 18.370 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1446.310 1685.620 1446.630 1685.680 ;
        RECT 1447.690 1685.620 1448.010 1685.680 ;
        RECT 1446.310 1685.480 1448.010 1685.620 ;
        RECT 1446.310 1685.420 1446.630 1685.480 ;
        RECT 1447.690 1685.420 1448.010 1685.480 ;
        RECT 1447.690 1659.440 1448.010 1659.500 ;
        RECT 2873.690 1659.440 2874.010 1659.500 ;
        RECT 1447.690 1659.300 2874.010 1659.440 ;
        RECT 1447.690 1659.240 1448.010 1659.300 ;
        RECT 2873.690 1659.240 2874.010 1659.300 ;
        RECT 2873.690 17.920 2874.010 17.980 ;
        RECT 2881.050 17.920 2881.370 17.980 ;
        RECT 2873.690 17.780 2881.370 17.920 ;
        RECT 2873.690 17.720 2874.010 17.780 ;
        RECT 2881.050 17.720 2881.370 17.780 ;
      LAYER via ;
        RECT 1446.340 1685.420 1446.600 1685.680 ;
        RECT 1447.720 1685.420 1447.980 1685.680 ;
        RECT 1447.720 1659.240 1447.980 1659.500 ;
        RECT 2873.720 1659.240 2873.980 1659.500 ;
        RECT 2873.720 17.720 2873.980 17.980 ;
        RECT 2881.080 17.720 2881.340 17.980 ;
      LAYER met2 ;
        RECT 1446.240 1700.340 1446.520 1704.000 ;
        RECT 1446.240 1700.000 1446.540 1700.340 ;
        RECT 1446.400 1685.710 1446.540 1700.000 ;
        RECT 1446.340 1685.390 1446.600 1685.710 ;
        RECT 1447.720 1685.390 1447.980 1685.710 ;
        RECT 1447.780 1659.530 1447.920 1685.390 ;
        RECT 1447.720 1659.210 1447.980 1659.530 ;
        RECT 2873.720 1659.210 2873.980 1659.530 ;
        RECT 2873.780 18.010 2873.920 1659.210 ;
        RECT 2873.720 17.690 2873.980 18.010 ;
        RECT 2881.080 17.690 2881.340 18.010 ;
        RECT 2881.140 2.400 2881.280 17.690 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1448.150 1673.040 1448.470 1673.100 ;
        RECT 2866.790 1673.040 2867.110 1673.100 ;
        RECT 1448.150 1672.900 2867.110 1673.040 ;
        RECT 1448.150 1672.840 1448.470 1672.900 ;
        RECT 2866.790 1672.840 2867.110 1672.900 ;
        RECT 2866.790 18.600 2867.110 18.660 ;
        RECT 2898.990 18.600 2899.310 18.660 ;
        RECT 2866.790 18.460 2899.310 18.600 ;
        RECT 2866.790 18.400 2867.110 18.460 ;
        RECT 2898.990 18.400 2899.310 18.460 ;
      LAYER via ;
        RECT 1448.180 1672.840 1448.440 1673.100 ;
        RECT 2866.820 1672.840 2867.080 1673.100 ;
        RECT 2866.820 18.400 2867.080 18.660 ;
        RECT 2899.020 18.400 2899.280 18.660 ;
      LAYER met2 ;
        RECT 1448.080 1700.340 1448.360 1704.000 ;
        RECT 1448.080 1700.000 1448.380 1700.340 ;
        RECT 1448.240 1673.130 1448.380 1700.000 ;
        RECT 1448.180 1672.810 1448.440 1673.130 ;
        RECT 2866.820 1672.810 2867.080 1673.130 ;
        RECT 2866.880 18.690 2867.020 1672.810 ;
        RECT 2866.820 18.370 2867.080 18.690 ;
        RECT 2899.020 18.370 2899.280 18.690 ;
        RECT 2899.080 2.400 2899.220 18.370 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 848.310 1681.200 848.630 1681.260 ;
        RECT 1236.550 1681.200 1236.870 1681.260 ;
        RECT 848.310 1681.060 1236.870 1681.200 ;
        RECT 848.310 1681.000 848.630 1681.060 ;
        RECT 1236.550 1681.000 1236.870 1681.060 ;
      LAYER via ;
        RECT 848.340 1681.000 848.600 1681.260 ;
        RECT 1236.580 1681.000 1236.840 1681.260 ;
      LAYER met2 ;
        RECT 1236.480 1700.340 1236.760 1704.000 ;
        RECT 1236.480 1700.000 1236.780 1700.340 ;
        RECT 1236.640 1681.290 1236.780 1700.000 ;
        RECT 848.340 1680.970 848.600 1681.290 ;
        RECT 1236.580 1680.970 1236.840 1681.290 ;
        RECT 848.400 17.410 848.540 1680.970 ;
        RECT 847.020 17.270 848.540 17.410 ;
        RECT 847.020 2.400 847.160 17.270 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1237.010 1691.060 1237.330 1691.120 ;
        RECT 1238.390 1691.060 1238.710 1691.120 ;
        RECT 1237.010 1690.920 1238.710 1691.060 ;
        RECT 1237.010 1690.860 1237.330 1690.920 ;
        RECT 1238.390 1690.860 1238.710 1690.920 ;
        RECT 1237.010 1668.080 1237.330 1668.340 ;
        RECT 869.010 1667.600 869.330 1667.660 ;
        RECT 1237.100 1667.600 1237.240 1668.080 ;
        RECT 869.010 1667.460 1237.240 1667.600 ;
        RECT 869.010 1667.400 869.330 1667.460 ;
      LAYER via ;
        RECT 1237.040 1690.860 1237.300 1691.120 ;
        RECT 1238.420 1690.860 1238.680 1691.120 ;
        RECT 1237.040 1668.080 1237.300 1668.340 ;
        RECT 869.040 1667.400 869.300 1667.660 ;
      LAYER met2 ;
        RECT 1238.320 1700.340 1238.600 1704.000 ;
        RECT 1238.320 1700.000 1238.620 1700.340 ;
        RECT 1238.480 1691.150 1238.620 1700.000 ;
        RECT 1237.040 1690.830 1237.300 1691.150 ;
        RECT 1238.420 1690.830 1238.680 1691.150 ;
        RECT 1237.100 1668.370 1237.240 1690.830 ;
        RECT 1237.040 1668.050 1237.300 1668.370 ;
        RECT 869.040 1667.370 869.300 1667.690 ;
        RECT 869.100 24.210 869.240 1667.370 ;
        RECT 864.960 24.070 869.240 24.210 ;
        RECT 864.960 2.400 865.100 24.070 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.810 1674.400 883.130 1674.460 ;
        RECT 1240.230 1674.400 1240.550 1674.460 ;
        RECT 882.810 1674.260 1240.550 1674.400 ;
        RECT 882.810 1674.200 883.130 1674.260 ;
        RECT 1240.230 1674.200 1240.550 1674.260 ;
      LAYER via ;
        RECT 882.840 1674.200 883.100 1674.460 ;
        RECT 1240.260 1674.200 1240.520 1674.460 ;
      LAYER met2 ;
        RECT 1240.160 1700.340 1240.440 1704.000 ;
        RECT 1240.160 1700.000 1240.460 1700.340 ;
        RECT 1240.320 1674.490 1240.460 1700.000 ;
        RECT 882.840 1674.170 883.100 1674.490 ;
        RECT 1240.260 1674.170 1240.520 1674.490 ;
        RECT 882.900 2.400 883.040 1674.170 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 903.510 1681.540 903.830 1681.600 ;
        RECT 1242.070 1681.540 1242.390 1681.600 ;
        RECT 903.510 1681.400 1242.390 1681.540 ;
        RECT 903.510 1681.340 903.830 1681.400 ;
        RECT 1242.070 1681.340 1242.390 1681.400 ;
      LAYER via ;
        RECT 903.540 1681.340 903.800 1681.600 ;
        RECT 1242.100 1681.340 1242.360 1681.600 ;
      LAYER met2 ;
        RECT 1242.000 1700.340 1242.280 1704.000 ;
        RECT 1242.000 1700.000 1242.300 1700.340 ;
        RECT 1242.160 1681.630 1242.300 1700.000 ;
        RECT 903.540 1681.310 903.800 1681.630 ;
        RECT 1242.100 1681.310 1242.360 1681.630 ;
        RECT 903.600 24.210 903.740 1681.310 ;
        RECT 900.840 24.070 903.740 24.210 ;
        RECT 900.840 2.400 900.980 24.070 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1243.985 1660.645 1244.155 1678.495 ;
      LAYER mcon ;
        RECT 1243.985 1678.325 1244.155 1678.495 ;
      LAYER met1 ;
        RECT 1243.910 1678.480 1244.230 1678.540 ;
        RECT 1243.715 1678.340 1244.230 1678.480 ;
        RECT 1243.910 1678.280 1244.230 1678.340 ;
        RECT 924.210 1660.800 924.530 1660.860 ;
        RECT 1243.925 1660.800 1244.215 1660.845 ;
        RECT 924.210 1660.660 1244.215 1660.800 ;
        RECT 924.210 1660.600 924.530 1660.660 ;
        RECT 1243.925 1660.615 1244.215 1660.660 ;
        RECT 918.690 2.960 919.010 3.020 ;
        RECT 923.750 2.960 924.070 3.020 ;
        RECT 918.690 2.820 924.070 2.960 ;
        RECT 918.690 2.760 919.010 2.820 ;
        RECT 923.750 2.760 924.070 2.820 ;
      LAYER via ;
        RECT 1243.940 1678.280 1244.200 1678.540 ;
        RECT 924.240 1660.600 924.500 1660.860 ;
        RECT 918.720 2.760 918.980 3.020 ;
        RECT 923.780 2.760 924.040 3.020 ;
      LAYER met2 ;
        RECT 1243.840 1700.340 1244.120 1704.000 ;
        RECT 1243.840 1700.000 1244.140 1700.340 ;
        RECT 1244.000 1678.570 1244.140 1700.000 ;
        RECT 1243.940 1678.250 1244.200 1678.570 ;
        RECT 924.240 1660.570 924.500 1660.890 ;
        RECT 924.300 33.730 924.440 1660.570 ;
        RECT 923.840 33.590 924.440 33.730 ;
        RECT 923.840 3.050 923.980 33.590 ;
        RECT 918.720 2.730 918.980 3.050 ;
        RECT 923.780 2.730 924.040 3.050 ;
        RECT 918.780 2.400 918.920 2.730 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1246.210 1678.140 1246.530 1678.200 ;
        RECT 1248.050 1678.140 1248.370 1678.200 ;
        RECT 1246.210 1678.000 1248.370 1678.140 ;
        RECT 1246.210 1677.940 1246.530 1678.000 ;
        RECT 1248.050 1677.940 1248.370 1678.000 ;
        RECT 936.170 26.420 936.490 26.480 ;
        RECT 1248.050 26.420 1248.370 26.480 ;
        RECT 936.170 26.280 1248.370 26.420 ;
        RECT 936.170 26.220 936.490 26.280 ;
        RECT 1248.050 26.220 1248.370 26.280 ;
      LAYER via ;
        RECT 1246.240 1677.940 1246.500 1678.200 ;
        RECT 1248.080 1677.940 1248.340 1678.200 ;
        RECT 936.200 26.220 936.460 26.480 ;
        RECT 1248.080 26.220 1248.340 26.480 ;
      LAYER met2 ;
        RECT 1245.680 1700.410 1245.960 1704.000 ;
        RECT 1245.680 1700.270 1246.440 1700.410 ;
        RECT 1245.680 1700.000 1245.960 1700.270 ;
        RECT 1246.300 1678.230 1246.440 1700.270 ;
        RECT 1246.240 1677.910 1246.500 1678.230 ;
        RECT 1248.080 1677.910 1248.340 1678.230 ;
        RECT 1248.140 26.510 1248.280 1677.910 ;
        RECT 936.200 26.190 936.460 26.510 ;
        RECT 1248.080 26.190 1248.340 26.510 ;
        RECT 936.260 2.400 936.400 26.190 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 954.110 26.760 954.430 26.820 ;
        RECT 1247.590 26.760 1247.910 26.820 ;
        RECT 954.110 26.620 1247.910 26.760 ;
        RECT 954.110 26.560 954.430 26.620 ;
        RECT 1247.590 26.560 1247.910 26.620 ;
      LAYER via ;
        RECT 954.140 26.560 954.400 26.820 ;
        RECT 1247.620 26.560 1247.880 26.820 ;
      LAYER met2 ;
        RECT 1247.520 1700.340 1247.800 1704.000 ;
        RECT 1247.520 1700.000 1247.820 1700.340 ;
        RECT 1247.680 26.850 1247.820 1700.000 ;
        RECT 954.140 26.530 954.400 26.850 ;
        RECT 1247.620 26.530 1247.880 26.850 ;
        RECT 954.200 2.400 954.340 26.530 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1221.445 25.925 1221.615 27.115 ;
      LAYER mcon ;
        RECT 1221.445 26.945 1221.615 27.115 ;
      LAYER met1 ;
        RECT 972.050 27.100 972.370 27.160 ;
        RECT 1221.385 27.100 1221.675 27.145 ;
        RECT 972.050 26.960 1221.675 27.100 ;
        RECT 972.050 26.900 972.370 26.960 ;
        RECT 1221.385 26.915 1221.675 26.960 ;
        RECT 1221.385 26.080 1221.675 26.125 ;
        RECT 1249.890 26.080 1250.210 26.140 ;
        RECT 1221.385 25.940 1250.210 26.080 ;
        RECT 1221.385 25.895 1221.675 25.940 ;
        RECT 1249.890 25.880 1250.210 25.940 ;
      LAYER via ;
        RECT 972.080 26.900 972.340 27.160 ;
        RECT 1249.920 25.880 1250.180 26.140 ;
      LAYER met2 ;
        RECT 1249.360 1700.410 1249.640 1704.000 ;
        RECT 1249.360 1700.270 1250.120 1700.410 ;
        RECT 1249.360 1700.000 1249.640 1700.270 ;
        RECT 972.080 26.870 972.340 27.190 ;
        RECT 972.140 2.400 972.280 26.870 ;
        RECT 1249.980 26.170 1250.120 1700.270 ;
        RECT 1249.920 25.850 1250.180 26.170 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 650.970 25.400 651.290 25.460 ;
        RECT 1217.230 25.400 1217.550 25.460 ;
        RECT 650.970 25.260 1217.550 25.400 ;
        RECT 650.970 25.200 651.290 25.260 ;
        RECT 1217.230 25.200 1217.550 25.260 ;
      LAYER via ;
        RECT 651.000 25.200 651.260 25.460 ;
        RECT 1217.260 25.200 1217.520 25.460 ;
      LAYER met2 ;
        RECT 1216.700 1700.340 1216.980 1704.000 ;
        RECT 1216.700 1700.000 1217.000 1700.340 ;
        RECT 1216.860 1677.290 1217.000 1700.000 ;
        RECT 1216.860 1677.150 1217.460 1677.290 ;
        RECT 1217.320 25.490 1217.460 1677.150 ;
        RECT 651.000 25.170 651.260 25.490 ;
        RECT 1217.260 25.170 1217.520 25.490 ;
        RECT 651.060 2.400 651.200 25.170 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1248.970 1677.460 1249.290 1677.520 ;
        RECT 1251.270 1677.460 1251.590 1677.520 ;
        RECT 1248.970 1677.320 1251.590 1677.460 ;
        RECT 1248.970 1677.260 1249.290 1677.320 ;
        RECT 1251.270 1677.260 1251.590 1677.320 ;
        RECT 989.990 27.440 990.310 27.500 ;
        RECT 989.990 27.300 1222.060 27.440 ;
        RECT 989.990 27.240 990.310 27.300 ;
        RECT 1221.920 27.100 1222.060 27.300 ;
        RECT 1248.970 27.100 1249.290 27.160 ;
        RECT 1221.920 26.960 1249.290 27.100 ;
        RECT 1248.970 26.900 1249.290 26.960 ;
      LAYER via ;
        RECT 1249.000 1677.260 1249.260 1677.520 ;
        RECT 1251.300 1677.260 1251.560 1677.520 ;
        RECT 990.020 27.240 990.280 27.500 ;
        RECT 1249.000 26.900 1249.260 27.160 ;
      LAYER met2 ;
        RECT 1251.200 1700.340 1251.480 1704.000 ;
        RECT 1251.200 1700.000 1251.500 1700.340 ;
        RECT 1251.360 1677.550 1251.500 1700.000 ;
        RECT 1249.000 1677.230 1249.260 1677.550 ;
        RECT 1251.300 1677.230 1251.560 1677.550 ;
        RECT 990.020 27.210 990.280 27.530 ;
        RECT 990.080 2.400 990.220 27.210 ;
        RECT 1249.060 27.190 1249.200 1677.230 ;
        RECT 1249.000 26.870 1249.260 27.190 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1255.485 351.985 1255.655 386.155 ;
      LAYER mcon ;
        RECT 1255.485 385.985 1255.655 386.155 ;
      LAYER met1 ;
        RECT 1253.570 1678.140 1253.890 1678.200 ;
        RECT 1255.410 1678.140 1255.730 1678.200 ;
        RECT 1253.570 1678.000 1255.730 1678.140 ;
        RECT 1253.570 1677.940 1253.890 1678.000 ;
        RECT 1255.410 1677.940 1255.730 1678.000 ;
        RECT 1255.410 386.140 1255.730 386.200 ;
        RECT 1255.215 386.000 1255.730 386.140 ;
        RECT 1255.410 385.940 1255.730 386.000 ;
        RECT 1255.410 352.140 1255.730 352.200 ;
        RECT 1255.215 352.000 1255.730 352.140 ;
        RECT 1255.410 351.940 1255.730 352.000 ;
        RECT 1007.470 23.700 1007.790 23.760 ;
        RECT 1255.410 23.700 1255.730 23.760 ;
        RECT 1007.470 23.560 1255.730 23.700 ;
        RECT 1007.470 23.500 1007.790 23.560 ;
        RECT 1255.410 23.500 1255.730 23.560 ;
      LAYER via ;
        RECT 1253.600 1677.940 1253.860 1678.200 ;
        RECT 1255.440 1677.940 1255.700 1678.200 ;
        RECT 1255.440 385.940 1255.700 386.200 ;
        RECT 1255.440 351.940 1255.700 352.200 ;
        RECT 1007.500 23.500 1007.760 23.760 ;
        RECT 1255.440 23.500 1255.700 23.760 ;
      LAYER met2 ;
        RECT 1253.040 1700.410 1253.320 1704.000 ;
        RECT 1253.040 1700.270 1253.800 1700.410 ;
        RECT 1253.040 1700.000 1253.320 1700.270 ;
        RECT 1253.660 1678.230 1253.800 1700.270 ;
        RECT 1253.600 1677.910 1253.860 1678.230 ;
        RECT 1255.440 1677.910 1255.700 1678.230 ;
        RECT 1255.500 386.230 1255.640 1677.910 ;
        RECT 1255.440 385.910 1255.700 386.230 ;
        RECT 1255.440 351.910 1255.700 352.230 ;
        RECT 1255.500 23.790 1255.640 351.910 ;
        RECT 1007.500 23.470 1007.760 23.790 ;
        RECT 1255.440 23.470 1255.700 23.790 ;
        RECT 1007.560 2.400 1007.700 23.470 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1255.025 358.445 1255.195 385.815 ;
      LAYER mcon ;
        RECT 1255.025 385.645 1255.195 385.815 ;
      LAYER met1 ;
        RECT 1254.950 385.800 1255.270 385.860 ;
        RECT 1254.755 385.660 1255.270 385.800 ;
        RECT 1254.950 385.600 1255.270 385.660 ;
        RECT 1254.950 358.600 1255.270 358.660 ;
        RECT 1254.755 358.460 1255.270 358.600 ;
        RECT 1254.950 358.400 1255.270 358.460 ;
        RECT 1025.410 23.360 1025.730 23.420 ;
        RECT 1254.950 23.360 1255.270 23.420 ;
        RECT 1025.410 23.220 1255.270 23.360 ;
        RECT 1025.410 23.160 1025.730 23.220 ;
        RECT 1254.950 23.160 1255.270 23.220 ;
      LAYER via ;
        RECT 1254.980 385.600 1255.240 385.860 ;
        RECT 1254.980 358.400 1255.240 358.660 ;
        RECT 1025.440 23.160 1025.700 23.420 ;
        RECT 1254.980 23.160 1255.240 23.420 ;
      LAYER met2 ;
        RECT 1254.880 1700.340 1255.160 1704.000 ;
        RECT 1254.880 1700.000 1255.180 1700.340 ;
        RECT 1255.040 385.890 1255.180 1700.000 ;
        RECT 1254.980 385.570 1255.240 385.890 ;
        RECT 1254.980 358.370 1255.240 358.690 ;
        RECT 1255.040 23.450 1255.180 358.370 ;
        RECT 1025.440 23.130 1025.700 23.450 ;
        RECT 1254.980 23.130 1255.240 23.450 ;
        RECT 1025.500 2.400 1025.640 23.130 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1214.470 1687.320 1214.790 1687.380 ;
        RECT 1256.790 1687.320 1257.110 1687.380 ;
        RECT 1214.470 1687.180 1257.110 1687.320 ;
        RECT 1214.470 1687.120 1214.790 1687.180 ;
        RECT 1256.790 1687.120 1257.110 1687.180 ;
        RECT 1048.410 1681.880 1048.730 1681.940 ;
        RECT 1214.470 1681.880 1214.790 1681.940 ;
        RECT 1048.410 1681.740 1214.790 1681.880 ;
        RECT 1048.410 1681.680 1048.730 1681.740 ;
        RECT 1214.470 1681.680 1214.790 1681.740 ;
        RECT 1043.350 2.960 1043.670 3.020 ;
        RECT 1048.410 2.960 1048.730 3.020 ;
        RECT 1043.350 2.820 1048.730 2.960 ;
        RECT 1043.350 2.760 1043.670 2.820 ;
        RECT 1048.410 2.760 1048.730 2.820 ;
      LAYER via ;
        RECT 1214.500 1687.120 1214.760 1687.380 ;
        RECT 1256.820 1687.120 1257.080 1687.380 ;
        RECT 1048.440 1681.680 1048.700 1681.940 ;
        RECT 1214.500 1681.680 1214.760 1681.940 ;
        RECT 1043.380 2.760 1043.640 3.020 ;
        RECT 1048.440 2.760 1048.700 3.020 ;
      LAYER met2 ;
        RECT 1256.720 1700.340 1257.000 1704.000 ;
        RECT 1256.720 1700.000 1257.020 1700.340 ;
        RECT 1256.880 1687.410 1257.020 1700.000 ;
        RECT 1214.500 1687.090 1214.760 1687.410 ;
        RECT 1256.820 1687.090 1257.080 1687.410 ;
        RECT 1214.560 1681.970 1214.700 1687.090 ;
        RECT 1048.440 1681.650 1048.700 1681.970 ;
        RECT 1214.500 1681.650 1214.760 1681.970 ;
        RECT 1048.500 3.050 1048.640 1681.650 ;
        RECT 1043.380 2.730 1043.640 3.050 ;
        RECT 1048.440 2.730 1048.700 3.050 ;
        RECT 1043.440 2.400 1043.580 2.730 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1258.705 1674.585 1258.875 1679.855 ;
      LAYER mcon ;
        RECT 1258.705 1679.685 1258.875 1679.855 ;
      LAYER met1 ;
        RECT 1258.630 1679.840 1258.950 1679.900 ;
        RECT 1258.435 1679.700 1258.950 1679.840 ;
        RECT 1258.630 1679.640 1258.950 1679.700 ;
        RECT 1062.210 1674.740 1062.530 1674.800 ;
        RECT 1258.645 1674.740 1258.935 1674.785 ;
        RECT 1062.210 1674.600 1258.935 1674.740 ;
        RECT 1062.210 1674.540 1062.530 1674.600 ;
        RECT 1258.645 1674.555 1258.935 1674.600 ;
      LAYER via ;
        RECT 1258.660 1679.640 1258.920 1679.900 ;
        RECT 1062.240 1674.540 1062.500 1674.800 ;
      LAYER met2 ;
        RECT 1258.560 1700.340 1258.840 1704.000 ;
        RECT 1258.560 1700.000 1258.860 1700.340 ;
        RECT 1258.720 1679.930 1258.860 1700.000 ;
        RECT 1258.660 1679.610 1258.920 1679.930 ;
        RECT 1062.240 1674.510 1062.500 1674.830 ;
        RECT 1062.300 18.090 1062.440 1674.510 ;
        RECT 1061.380 17.950 1062.440 18.090 ;
        RECT 1061.380 2.400 1061.520 17.950 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1260.930 1684.940 1261.250 1685.000 ;
        RECT 1262.770 1684.940 1263.090 1685.000 ;
        RECT 1260.930 1684.800 1263.090 1684.940 ;
        RECT 1260.930 1684.740 1261.250 1684.800 ;
        RECT 1262.770 1684.740 1263.090 1684.800 ;
        RECT 1262.310 1668.620 1262.630 1668.680 ;
        RECT 1236.640 1668.480 1262.630 1668.620 ;
        RECT 1082.910 1667.940 1083.230 1668.000 ;
        RECT 1236.640 1667.940 1236.780 1668.480 ;
        RECT 1262.310 1668.420 1262.630 1668.480 ;
        RECT 1082.910 1667.800 1236.780 1667.940 ;
        RECT 1082.910 1667.740 1083.230 1667.800 ;
      LAYER via ;
        RECT 1260.960 1684.740 1261.220 1685.000 ;
        RECT 1262.800 1684.740 1263.060 1685.000 ;
        RECT 1082.940 1667.740 1083.200 1668.000 ;
        RECT 1262.340 1668.420 1262.600 1668.680 ;
      LAYER met2 ;
        RECT 1260.400 1700.410 1260.680 1704.000 ;
        RECT 1260.400 1700.270 1261.160 1700.410 ;
        RECT 1260.400 1700.000 1260.680 1700.270 ;
        RECT 1261.020 1685.030 1261.160 1700.270 ;
        RECT 1260.960 1684.710 1261.220 1685.030 ;
        RECT 1262.800 1684.710 1263.060 1685.030 ;
        RECT 1262.860 1681.370 1263.000 1684.710 ;
        RECT 1262.400 1681.230 1263.000 1681.370 ;
        RECT 1262.400 1668.710 1262.540 1681.230 ;
        RECT 1262.340 1668.390 1262.600 1668.710 ;
        RECT 1082.940 1667.710 1083.200 1668.030 ;
        RECT 1083.000 18.090 1083.140 1667.710 ;
        RECT 1079.320 17.950 1083.140 18.090 ;
        RECT 1079.320 2.400 1079.460 17.950 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1096.710 1682.220 1097.030 1682.280 ;
        RECT 1262.310 1682.220 1262.630 1682.280 ;
        RECT 1096.710 1682.080 1262.630 1682.220 ;
        RECT 1096.710 1682.020 1097.030 1682.080 ;
        RECT 1262.310 1682.020 1262.630 1682.080 ;
      LAYER via ;
        RECT 1096.740 1682.020 1097.000 1682.280 ;
        RECT 1262.340 1682.020 1262.600 1682.280 ;
      LAYER met2 ;
        RECT 1262.240 1700.340 1262.520 1704.000 ;
        RECT 1262.240 1700.000 1262.540 1700.340 ;
        RECT 1262.400 1682.310 1262.540 1700.000 ;
        RECT 1096.740 1681.990 1097.000 1682.310 ;
        RECT 1262.340 1681.990 1262.600 1682.310 ;
        RECT 1096.800 2.400 1096.940 1681.990 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1117.410 1675.080 1117.730 1675.140 ;
        RECT 1264.150 1675.080 1264.470 1675.140 ;
        RECT 1117.410 1674.940 1264.470 1675.080 ;
        RECT 1117.410 1674.880 1117.730 1674.940 ;
        RECT 1264.150 1674.880 1264.470 1674.940 ;
      LAYER via ;
        RECT 1117.440 1674.880 1117.700 1675.140 ;
        RECT 1264.180 1674.880 1264.440 1675.140 ;
      LAYER met2 ;
        RECT 1264.080 1700.340 1264.360 1704.000 ;
        RECT 1264.080 1700.000 1264.380 1700.340 ;
        RECT 1264.240 1675.170 1264.380 1700.000 ;
        RECT 1117.440 1674.850 1117.700 1675.170 ;
        RECT 1264.180 1674.850 1264.440 1675.170 ;
        RECT 1117.500 16.730 1117.640 1674.850 ;
        RECT 1114.740 16.590 1117.640 16.730 ;
        RECT 1114.740 2.400 1114.880 16.590 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1265.070 1690.720 1265.390 1690.780 ;
        RECT 1265.990 1690.720 1266.310 1690.780 ;
        RECT 1265.070 1690.580 1266.310 1690.720 ;
        RECT 1265.070 1690.520 1265.390 1690.580 ;
        RECT 1265.990 1690.520 1266.310 1690.580 ;
        RECT 1159.730 1686.980 1160.050 1687.040 ;
        RECT 1265.070 1686.980 1265.390 1687.040 ;
        RECT 1159.730 1686.840 1265.390 1686.980 ;
        RECT 1159.730 1686.780 1160.050 1686.840 ;
        RECT 1265.070 1686.780 1265.390 1686.840 ;
        RECT 1138.110 1676.780 1138.430 1676.840 ;
        RECT 1159.730 1676.780 1160.050 1676.840 ;
        RECT 1138.110 1676.640 1160.050 1676.780 ;
        RECT 1138.110 1676.580 1138.430 1676.640 ;
        RECT 1159.730 1676.580 1160.050 1676.640 ;
        RECT 1132.590 19.280 1132.910 19.340 ;
        RECT 1138.110 19.280 1138.430 19.340 ;
        RECT 1132.590 19.140 1138.430 19.280 ;
        RECT 1132.590 19.080 1132.910 19.140 ;
        RECT 1138.110 19.080 1138.430 19.140 ;
      LAYER via ;
        RECT 1265.100 1690.520 1265.360 1690.780 ;
        RECT 1266.020 1690.520 1266.280 1690.780 ;
        RECT 1159.760 1686.780 1160.020 1687.040 ;
        RECT 1265.100 1686.780 1265.360 1687.040 ;
        RECT 1138.140 1676.580 1138.400 1676.840 ;
        RECT 1159.760 1676.580 1160.020 1676.840 ;
        RECT 1132.620 19.080 1132.880 19.340 ;
        RECT 1138.140 19.080 1138.400 19.340 ;
      LAYER met2 ;
        RECT 1265.920 1700.340 1266.200 1704.000 ;
        RECT 1265.920 1700.000 1266.220 1700.340 ;
        RECT 1266.080 1690.810 1266.220 1700.000 ;
        RECT 1265.100 1690.490 1265.360 1690.810 ;
        RECT 1266.020 1690.490 1266.280 1690.810 ;
        RECT 1265.160 1687.070 1265.300 1690.490 ;
        RECT 1159.760 1686.750 1160.020 1687.070 ;
        RECT 1265.100 1686.750 1265.360 1687.070 ;
        RECT 1159.820 1676.870 1159.960 1686.750 ;
        RECT 1138.140 1676.550 1138.400 1676.870 ;
        RECT 1159.760 1676.550 1160.020 1676.870 ;
        RECT 1138.200 19.370 1138.340 1676.550 ;
        RECT 1132.620 19.050 1132.880 19.370 ;
        RECT 1138.140 19.050 1138.400 19.370 ;
        RECT 1132.680 2.400 1132.820 19.050 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1152.370 1682.560 1152.690 1682.620 ;
        RECT 1267.830 1682.560 1268.150 1682.620 ;
        RECT 1152.370 1682.420 1268.150 1682.560 ;
        RECT 1152.370 1682.360 1152.690 1682.420 ;
        RECT 1267.830 1682.360 1268.150 1682.420 ;
        RECT 1150.530 2.960 1150.850 3.020 ;
        RECT 1151.910 2.960 1152.230 3.020 ;
        RECT 1150.530 2.820 1152.230 2.960 ;
        RECT 1150.530 2.760 1150.850 2.820 ;
        RECT 1151.910 2.760 1152.230 2.820 ;
      LAYER via ;
        RECT 1152.400 1682.360 1152.660 1682.620 ;
        RECT 1267.860 1682.360 1268.120 1682.620 ;
        RECT 1150.560 2.760 1150.820 3.020 ;
        RECT 1151.940 2.760 1152.200 3.020 ;
      LAYER met2 ;
        RECT 1267.760 1700.340 1268.040 1704.000 ;
        RECT 1267.760 1700.000 1268.060 1700.340 ;
        RECT 1267.920 1682.650 1268.060 1700.000 ;
        RECT 1152.400 1682.330 1152.660 1682.650 ;
        RECT 1267.860 1682.330 1268.120 1682.650 ;
        RECT 1152.460 1675.930 1152.600 1682.330 ;
        RECT 1152.000 1675.790 1152.600 1675.930 ;
        RECT 1152.000 3.050 1152.140 1675.790 ;
        RECT 1150.560 2.730 1150.820 3.050 ;
        RECT 1151.940 2.730 1152.200 3.050 ;
        RECT 1150.620 2.400 1150.760 2.730 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.910 25.740 669.230 25.800 ;
        RECT 1218.610 25.740 1218.930 25.800 ;
        RECT 668.910 25.600 1218.930 25.740 ;
        RECT 668.910 25.540 669.230 25.600 ;
        RECT 1218.610 25.540 1218.930 25.600 ;
      LAYER via ;
        RECT 668.940 25.540 669.200 25.800 ;
        RECT 1218.640 25.540 1218.900 25.800 ;
      LAYER met2 ;
        RECT 1218.540 1700.340 1218.820 1704.000 ;
        RECT 1218.540 1700.000 1218.840 1700.340 ;
        RECT 1218.700 25.830 1218.840 1700.000 ;
        RECT 668.940 25.510 669.200 25.830 ;
        RECT 1218.640 25.510 1218.900 25.830 ;
        RECT 669.000 2.400 669.140 25.510 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1270.130 1667.600 1270.450 1667.660 ;
        RECT 1271.050 1667.600 1271.370 1667.660 ;
        RECT 1270.130 1667.460 1271.370 1667.600 ;
        RECT 1270.130 1667.400 1270.450 1667.460 ;
        RECT 1271.050 1667.400 1271.370 1667.460 ;
        RECT 1168.470 24.040 1168.790 24.100 ;
        RECT 1271.050 24.040 1271.370 24.100 ;
        RECT 1168.470 23.900 1271.370 24.040 ;
        RECT 1168.470 23.840 1168.790 23.900 ;
        RECT 1271.050 23.840 1271.370 23.900 ;
      LAYER via ;
        RECT 1270.160 1667.400 1270.420 1667.660 ;
        RECT 1271.080 1667.400 1271.340 1667.660 ;
        RECT 1168.500 23.840 1168.760 24.100 ;
        RECT 1271.080 23.840 1271.340 24.100 ;
      LAYER met2 ;
        RECT 1269.600 1700.410 1269.880 1704.000 ;
        RECT 1269.600 1700.270 1270.360 1700.410 ;
        RECT 1269.600 1700.000 1269.880 1700.270 ;
        RECT 1270.220 1667.690 1270.360 1700.270 ;
        RECT 1270.160 1667.370 1270.420 1667.690 ;
        RECT 1271.080 1667.370 1271.340 1667.690 ;
        RECT 1271.140 24.130 1271.280 1667.370 ;
        RECT 1168.500 23.810 1168.760 24.130 ;
        RECT 1271.080 23.810 1271.340 24.130 ;
        RECT 1168.560 2.400 1168.700 23.810 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 24.380 1186.730 24.440 ;
        RECT 1270.590 24.380 1270.910 24.440 ;
        RECT 1186.410 24.240 1270.910 24.380 ;
        RECT 1186.410 24.180 1186.730 24.240 ;
        RECT 1270.590 24.180 1270.910 24.240 ;
      LAYER via ;
        RECT 1186.440 24.180 1186.700 24.440 ;
        RECT 1270.620 24.180 1270.880 24.440 ;
      LAYER met2 ;
        RECT 1271.440 1700.340 1271.720 1704.000 ;
        RECT 1271.440 1700.000 1271.740 1700.340 ;
        RECT 1271.600 1678.650 1271.740 1700.000 ;
        RECT 1270.680 1678.510 1271.740 1678.650 ;
        RECT 1270.680 24.470 1270.820 1678.510 ;
        RECT 1186.440 24.150 1186.700 24.470 ;
        RECT 1270.620 24.150 1270.880 24.470 ;
        RECT 1186.500 12.650 1186.640 24.150 ;
        RECT 1186.040 12.510 1186.640 12.650 ;
        RECT 1186.040 2.400 1186.180 12.510 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1271.510 1678.140 1271.830 1678.200 ;
        RECT 1273.350 1678.140 1273.670 1678.200 ;
        RECT 1271.510 1678.000 1273.670 1678.140 ;
        RECT 1271.510 1677.940 1271.830 1678.000 ;
        RECT 1273.350 1677.940 1273.670 1678.000 ;
        RECT 1203.890 24.720 1204.210 24.780 ;
        RECT 1271.510 24.720 1271.830 24.780 ;
        RECT 1203.890 24.580 1271.830 24.720 ;
        RECT 1203.890 24.520 1204.210 24.580 ;
        RECT 1271.510 24.520 1271.830 24.580 ;
      LAYER via ;
        RECT 1271.540 1677.940 1271.800 1678.200 ;
        RECT 1273.380 1677.940 1273.640 1678.200 ;
        RECT 1203.920 24.520 1204.180 24.780 ;
        RECT 1271.540 24.520 1271.800 24.780 ;
      LAYER met2 ;
        RECT 1273.280 1700.340 1273.560 1704.000 ;
        RECT 1273.280 1700.000 1273.580 1700.340 ;
        RECT 1273.440 1678.230 1273.580 1700.000 ;
        RECT 1271.540 1677.910 1271.800 1678.230 ;
        RECT 1273.380 1677.910 1273.640 1678.230 ;
        RECT 1271.600 24.810 1271.740 1677.910 ;
        RECT 1203.920 24.490 1204.180 24.810 ;
        RECT 1271.540 24.490 1271.800 24.810 ;
        RECT 1203.980 2.400 1204.120 24.490 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1238.390 1690.380 1238.710 1690.440 ;
        RECT 1275.190 1690.380 1275.510 1690.440 ;
        RECT 1238.390 1690.240 1275.510 1690.380 ;
        RECT 1238.390 1690.180 1238.710 1690.240 ;
        RECT 1275.190 1690.180 1275.510 1690.240 ;
        RECT 1221.830 25.740 1222.150 25.800 ;
        RECT 1238.390 25.740 1238.710 25.800 ;
        RECT 1221.830 25.600 1238.710 25.740 ;
        RECT 1221.830 25.540 1222.150 25.600 ;
        RECT 1238.390 25.540 1238.710 25.600 ;
      LAYER via ;
        RECT 1238.420 1690.180 1238.680 1690.440 ;
        RECT 1275.220 1690.180 1275.480 1690.440 ;
        RECT 1221.860 25.540 1222.120 25.800 ;
        RECT 1238.420 25.540 1238.680 25.800 ;
      LAYER met2 ;
        RECT 1275.120 1700.340 1275.400 1704.000 ;
        RECT 1275.120 1700.000 1275.420 1700.340 ;
        RECT 1275.280 1690.470 1275.420 1700.000 ;
        RECT 1238.420 1690.150 1238.680 1690.470 ;
        RECT 1275.220 1690.150 1275.480 1690.470 ;
        RECT 1238.480 25.830 1238.620 1690.150 ;
        RECT 1221.860 25.510 1222.120 25.830 ;
        RECT 1238.420 25.510 1238.680 25.830 ;
        RECT 1221.920 2.400 1222.060 25.510 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1272.890 1683.920 1273.210 1683.980 ;
        RECT 1277.030 1683.920 1277.350 1683.980 ;
        RECT 1272.890 1683.780 1277.350 1683.920 ;
        RECT 1272.890 1683.720 1273.210 1683.780 ;
        RECT 1277.030 1683.720 1277.350 1683.780 ;
        RECT 1239.770 18.260 1240.090 18.320 ;
        RECT 1272.890 18.260 1273.210 18.320 ;
        RECT 1239.770 18.120 1273.210 18.260 ;
        RECT 1239.770 18.060 1240.090 18.120 ;
        RECT 1272.890 18.060 1273.210 18.120 ;
      LAYER via ;
        RECT 1272.920 1683.720 1273.180 1683.980 ;
        RECT 1277.060 1683.720 1277.320 1683.980 ;
        RECT 1239.800 18.060 1240.060 18.320 ;
        RECT 1272.920 18.060 1273.180 18.320 ;
      LAYER met2 ;
        RECT 1276.960 1700.340 1277.240 1704.000 ;
        RECT 1276.960 1700.000 1277.260 1700.340 ;
        RECT 1277.120 1684.010 1277.260 1700.000 ;
        RECT 1272.920 1683.690 1273.180 1684.010 ;
        RECT 1277.060 1683.690 1277.320 1684.010 ;
        RECT 1272.980 18.350 1273.120 1683.690 ;
        RECT 1239.800 18.030 1240.060 18.350 ;
        RECT 1272.920 18.030 1273.180 18.350 ;
        RECT 1239.860 2.400 1240.000 18.030 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1273.425 1642.285 1273.595 1678.835 ;
      LAYER mcon ;
        RECT 1273.425 1678.665 1273.595 1678.835 ;
      LAYER met1 ;
        RECT 1273.365 1678.820 1273.655 1678.865 ;
        RECT 1278.870 1678.820 1279.190 1678.880 ;
        RECT 1273.365 1678.680 1279.190 1678.820 ;
        RECT 1273.365 1678.635 1273.655 1678.680 ;
        RECT 1278.870 1678.620 1279.190 1678.680 ;
        RECT 1273.350 1642.440 1273.670 1642.500 ;
        RECT 1273.155 1642.300 1273.670 1642.440 ;
        RECT 1273.350 1642.240 1273.670 1642.300 ;
        RECT 1257.250 2.960 1257.570 3.020 ;
        RECT 1273.350 2.960 1273.670 3.020 ;
        RECT 1257.250 2.820 1273.670 2.960 ;
        RECT 1257.250 2.760 1257.570 2.820 ;
        RECT 1273.350 2.760 1273.670 2.820 ;
      LAYER via ;
        RECT 1278.900 1678.620 1279.160 1678.880 ;
        RECT 1273.380 1642.240 1273.640 1642.500 ;
        RECT 1257.280 2.760 1257.540 3.020 ;
        RECT 1273.380 2.760 1273.640 3.020 ;
      LAYER met2 ;
        RECT 1278.800 1700.340 1279.080 1704.000 ;
        RECT 1278.800 1700.000 1279.100 1700.340 ;
        RECT 1278.960 1678.910 1279.100 1700.000 ;
        RECT 1278.900 1678.590 1279.160 1678.910 ;
        RECT 1273.380 1642.210 1273.640 1642.530 ;
        RECT 1273.440 3.050 1273.580 1642.210 ;
        RECT 1257.280 2.730 1257.540 3.050 ;
        RECT 1273.380 2.730 1273.640 3.050 ;
        RECT 1257.340 2.400 1257.480 2.730 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1275.190 20.640 1275.510 20.700 ;
        RECT 1280.710 20.640 1281.030 20.700 ;
        RECT 1275.190 20.500 1281.030 20.640 ;
        RECT 1275.190 20.440 1275.510 20.500 ;
        RECT 1280.710 20.440 1281.030 20.500 ;
      LAYER via ;
        RECT 1275.220 20.440 1275.480 20.700 ;
        RECT 1280.740 20.440 1281.000 20.700 ;
      LAYER met2 ;
        RECT 1280.640 1700.340 1280.920 1704.000 ;
        RECT 1280.640 1700.000 1280.940 1700.340 ;
        RECT 1280.800 20.730 1280.940 1700.000 ;
        RECT 1275.220 20.410 1275.480 20.730 ;
        RECT 1280.740 20.410 1281.000 20.730 ;
        RECT 1275.280 2.400 1275.420 20.410 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1282.550 1684.260 1282.870 1684.320 ;
        RECT 1286.690 1684.260 1287.010 1684.320 ;
        RECT 1282.550 1684.120 1287.010 1684.260 ;
        RECT 1282.550 1684.060 1282.870 1684.120 ;
        RECT 1286.690 1684.060 1287.010 1684.120 ;
        RECT 1286.690 20.300 1287.010 20.360 ;
        RECT 1293.130 20.300 1293.450 20.360 ;
        RECT 1286.690 20.160 1293.450 20.300 ;
        RECT 1286.690 20.100 1287.010 20.160 ;
        RECT 1293.130 20.100 1293.450 20.160 ;
      LAYER via ;
        RECT 1282.580 1684.060 1282.840 1684.320 ;
        RECT 1286.720 1684.060 1286.980 1684.320 ;
        RECT 1286.720 20.100 1286.980 20.360 ;
        RECT 1293.160 20.100 1293.420 20.360 ;
      LAYER met2 ;
        RECT 1282.480 1700.340 1282.760 1704.000 ;
        RECT 1282.480 1700.000 1282.780 1700.340 ;
        RECT 1282.640 1684.350 1282.780 1700.000 ;
        RECT 1282.580 1684.030 1282.840 1684.350 ;
        RECT 1286.720 1684.030 1286.980 1684.350 ;
        RECT 1286.780 20.390 1286.920 1684.030 ;
        RECT 1286.720 20.070 1286.980 20.390 ;
        RECT 1293.160 20.070 1293.420 20.390 ;
        RECT 1293.220 2.400 1293.360 20.070 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1286.305 572.645 1286.475 620.755 ;
        RECT 1286.305 469.285 1286.475 476.255 ;
        RECT 1285.845 317.645 1286.015 341.955 ;
        RECT 1285.845 172.465 1286.015 196.775 ;
        RECT 1286.305 89.845 1286.475 137.955 ;
      LAYER mcon ;
        RECT 1286.305 620.585 1286.475 620.755 ;
        RECT 1286.305 476.085 1286.475 476.255 ;
        RECT 1285.845 341.785 1286.015 341.955 ;
        RECT 1285.845 196.605 1286.015 196.775 ;
        RECT 1286.305 137.785 1286.475 137.955 ;
      LAYER met1 ;
        RECT 1284.390 1673.380 1284.710 1673.440 ;
        RECT 1285.770 1673.380 1286.090 1673.440 ;
        RECT 1284.390 1673.240 1286.090 1673.380 ;
        RECT 1284.390 1673.180 1284.710 1673.240 ;
        RECT 1285.770 1673.180 1286.090 1673.240 ;
        RECT 1285.770 1642.100 1286.090 1642.160 ;
        RECT 1286.230 1642.100 1286.550 1642.160 ;
        RECT 1285.770 1641.960 1286.550 1642.100 ;
        RECT 1285.770 1641.900 1286.090 1641.960 ;
        RECT 1286.230 1641.900 1286.550 1641.960 ;
        RECT 1285.770 1435.380 1286.090 1435.440 ;
        RECT 1286.230 1435.380 1286.550 1435.440 ;
        RECT 1285.770 1435.240 1286.550 1435.380 ;
        RECT 1285.770 1435.180 1286.090 1435.240 ;
        RECT 1286.230 1435.180 1286.550 1435.240 ;
        RECT 1285.770 1304.480 1286.090 1304.540 ;
        RECT 1286.230 1304.480 1286.550 1304.540 ;
        RECT 1285.770 1304.340 1286.550 1304.480 ;
        RECT 1285.770 1304.280 1286.090 1304.340 ;
        RECT 1286.230 1304.280 1286.550 1304.340 ;
        RECT 1284.850 1249.060 1285.170 1249.120 ;
        RECT 1286.230 1249.060 1286.550 1249.120 ;
        RECT 1284.850 1248.920 1286.550 1249.060 ;
        RECT 1284.850 1248.860 1285.170 1248.920 ;
        RECT 1286.230 1248.860 1286.550 1248.920 ;
        RECT 1286.230 845.480 1286.550 845.540 ;
        RECT 1287.150 845.480 1287.470 845.540 ;
        RECT 1286.230 845.340 1287.470 845.480 ;
        RECT 1286.230 845.280 1286.550 845.340 ;
        RECT 1287.150 845.280 1287.470 845.340 ;
        RECT 1286.230 773.400 1286.550 773.460 ;
        RECT 1285.860 773.260 1286.550 773.400 ;
        RECT 1285.860 772.780 1286.000 773.260 ;
        RECT 1286.230 773.200 1286.550 773.260 ;
        RECT 1285.770 772.520 1286.090 772.780 ;
        RECT 1285.770 651.820 1286.090 652.080 ;
        RECT 1285.860 651.680 1286.000 651.820 ;
        RECT 1286.230 651.680 1286.550 651.740 ;
        RECT 1285.860 651.540 1286.550 651.680 ;
        RECT 1286.230 651.480 1286.550 651.540 ;
        RECT 1286.230 620.740 1286.550 620.800 ;
        RECT 1286.035 620.600 1286.550 620.740 ;
        RECT 1286.230 620.540 1286.550 620.600 ;
        RECT 1286.230 572.800 1286.550 572.860 ;
        RECT 1286.035 572.660 1286.550 572.800 ;
        RECT 1286.230 572.600 1286.550 572.660 ;
        RECT 1286.230 476.240 1286.550 476.300 ;
        RECT 1286.035 476.100 1286.550 476.240 ;
        RECT 1286.230 476.040 1286.550 476.100 ;
        RECT 1286.230 469.440 1286.550 469.500 ;
        RECT 1286.035 469.300 1286.550 469.440 ;
        RECT 1286.230 469.240 1286.550 469.300 ;
        RECT 1285.785 341.940 1286.075 341.985 ;
        RECT 1286.230 341.940 1286.550 342.000 ;
        RECT 1285.785 341.800 1286.550 341.940 ;
        RECT 1285.785 341.755 1286.075 341.800 ;
        RECT 1286.230 341.740 1286.550 341.800 ;
        RECT 1285.770 317.800 1286.090 317.860 ;
        RECT 1285.575 317.660 1286.090 317.800 ;
        RECT 1285.770 317.600 1286.090 317.660 ;
        RECT 1284.850 262.380 1285.170 262.440 ;
        RECT 1286.230 262.380 1286.550 262.440 ;
        RECT 1284.850 262.240 1286.550 262.380 ;
        RECT 1284.850 262.180 1285.170 262.240 ;
        RECT 1286.230 262.180 1286.550 262.240 ;
        RECT 1285.770 241.640 1286.090 241.700 ;
        RECT 1286.230 241.640 1286.550 241.700 ;
        RECT 1285.770 241.500 1286.550 241.640 ;
        RECT 1285.770 241.440 1286.090 241.500 ;
        RECT 1286.230 241.440 1286.550 241.500 ;
        RECT 1285.770 196.760 1286.090 196.820 ;
        RECT 1285.575 196.620 1286.090 196.760 ;
        RECT 1285.770 196.560 1286.090 196.620 ;
        RECT 1285.785 172.620 1286.075 172.665 ;
        RECT 1286.230 172.620 1286.550 172.680 ;
        RECT 1285.785 172.480 1286.550 172.620 ;
        RECT 1285.785 172.435 1286.075 172.480 ;
        RECT 1286.230 172.420 1286.550 172.480 ;
        RECT 1286.230 137.940 1286.550 138.000 ;
        RECT 1286.035 137.800 1286.550 137.940 ;
        RECT 1286.230 137.740 1286.550 137.800 ;
        RECT 1286.230 90.000 1286.550 90.060 ;
        RECT 1286.035 89.860 1286.550 90.000 ;
        RECT 1286.230 89.800 1286.550 89.860 ;
        RECT 1285.770 48.520 1286.090 48.580 ;
        RECT 1286.230 48.520 1286.550 48.580 ;
        RECT 1285.770 48.380 1286.550 48.520 ;
        RECT 1285.770 48.320 1286.090 48.380 ;
        RECT 1286.230 48.320 1286.550 48.380 ;
        RECT 1285.770 19.620 1286.090 19.680 ;
        RECT 1311.070 19.620 1311.390 19.680 ;
        RECT 1285.770 19.480 1311.390 19.620 ;
        RECT 1285.770 19.420 1286.090 19.480 ;
        RECT 1311.070 19.420 1311.390 19.480 ;
      LAYER via ;
        RECT 1284.420 1673.180 1284.680 1673.440 ;
        RECT 1285.800 1673.180 1286.060 1673.440 ;
        RECT 1285.800 1641.900 1286.060 1642.160 ;
        RECT 1286.260 1641.900 1286.520 1642.160 ;
        RECT 1285.800 1435.180 1286.060 1435.440 ;
        RECT 1286.260 1435.180 1286.520 1435.440 ;
        RECT 1285.800 1304.280 1286.060 1304.540 ;
        RECT 1286.260 1304.280 1286.520 1304.540 ;
        RECT 1284.880 1248.860 1285.140 1249.120 ;
        RECT 1286.260 1248.860 1286.520 1249.120 ;
        RECT 1286.260 845.280 1286.520 845.540 ;
        RECT 1287.180 845.280 1287.440 845.540 ;
        RECT 1286.260 773.200 1286.520 773.460 ;
        RECT 1285.800 772.520 1286.060 772.780 ;
        RECT 1285.800 651.820 1286.060 652.080 ;
        RECT 1286.260 651.480 1286.520 651.740 ;
        RECT 1286.260 620.540 1286.520 620.800 ;
        RECT 1286.260 572.600 1286.520 572.860 ;
        RECT 1286.260 476.040 1286.520 476.300 ;
        RECT 1286.260 469.240 1286.520 469.500 ;
        RECT 1286.260 341.740 1286.520 342.000 ;
        RECT 1285.800 317.600 1286.060 317.860 ;
        RECT 1284.880 262.180 1285.140 262.440 ;
        RECT 1286.260 262.180 1286.520 262.440 ;
        RECT 1285.800 241.440 1286.060 241.700 ;
        RECT 1286.260 241.440 1286.520 241.700 ;
        RECT 1285.800 196.560 1286.060 196.820 ;
        RECT 1286.260 172.420 1286.520 172.680 ;
        RECT 1286.260 137.740 1286.520 138.000 ;
        RECT 1286.260 89.800 1286.520 90.060 ;
        RECT 1285.800 48.320 1286.060 48.580 ;
        RECT 1286.260 48.320 1286.520 48.580 ;
        RECT 1285.800 19.420 1286.060 19.680 ;
        RECT 1311.100 19.420 1311.360 19.680 ;
      LAYER met2 ;
        RECT 1284.320 1700.340 1284.600 1704.000 ;
        RECT 1284.320 1700.000 1284.620 1700.340 ;
        RECT 1284.480 1673.470 1284.620 1700.000 ;
        RECT 1284.420 1673.150 1284.680 1673.470 ;
        RECT 1285.800 1673.150 1286.060 1673.470 ;
        RECT 1285.860 1642.190 1286.000 1673.150 ;
        RECT 1285.800 1641.870 1286.060 1642.190 ;
        RECT 1286.260 1641.870 1286.520 1642.190 ;
        RECT 1286.320 1435.470 1286.460 1641.870 ;
        RECT 1285.800 1435.150 1286.060 1435.470 ;
        RECT 1286.260 1435.150 1286.520 1435.470 ;
        RECT 1285.860 1331.850 1286.000 1435.150 ;
        RECT 1285.860 1331.710 1286.460 1331.850 ;
        RECT 1286.320 1304.570 1286.460 1331.710 ;
        RECT 1285.800 1304.250 1286.060 1304.570 ;
        RECT 1286.260 1304.250 1286.520 1304.570 ;
        RECT 1285.860 1297.285 1286.000 1304.250 ;
        RECT 1284.870 1296.915 1285.150 1297.285 ;
        RECT 1285.790 1296.915 1286.070 1297.285 ;
        RECT 1284.940 1249.150 1285.080 1296.915 ;
        RECT 1284.880 1248.830 1285.140 1249.150 ;
        RECT 1286.260 1248.830 1286.520 1249.150 ;
        RECT 1286.320 1145.645 1286.460 1248.830 ;
        RECT 1286.250 1145.275 1286.530 1145.645 ;
        RECT 1286.250 1144.595 1286.530 1144.965 ;
        RECT 1286.320 845.570 1286.460 1144.595 ;
        RECT 1286.260 845.250 1286.520 845.570 ;
        RECT 1287.180 845.250 1287.440 845.570 ;
        RECT 1287.240 821.285 1287.380 845.250 ;
        RECT 1286.250 820.915 1286.530 821.285 ;
        RECT 1287.170 820.915 1287.450 821.285 ;
        RECT 1286.320 773.490 1286.460 820.915 ;
        RECT 1286.260 773.170 1286.520 773.490 ;
        RECT 1285.800 772.490 1286.060 772.810 ;
        RECT 1285.860 652.110 1286.000 772.490 ;
        RECT 1285.800 651.790 1286.060 652.110 ;
        RECT 1286.260 651.450 1286.520 651.770 ;
        RECT 1286.320 620.830 1286.460 651.450 ;
        RECT 1286.260 620.510 1286.520 620.830 ;
        RECT 1286.260 572.570 1286.520 572.890 ;
        RECT 1286.320 476.330 1286.460 572.570 ;
        RECT 1286.260 476.010 1286.520 476.330 ;
        RECT 1286.260 469.210 1286.520 469.530 ;
        RECT 1286.320 421.330 1286.460 469.210 ;
        RECT 1285.860 421.190 1286.460 421.330 ;
        RECT 1285.860 389.370 1286.000 421.190 ;
        RECT 1285.860 389.230 1286.460 389.370 ;
        RECT 1286.320 342.030 1286.460 389.230 ;
        RECT 1286.260 341.710 1286.520 342.030 ;
        RECT 1285.800 317.570 1286.060 317.890 ;
        RECT 1285.860 310.605 1286.000 317.570 ;
        RECT 1284.870 310.235 1285.150 310.605 ;
        RECT 1285.790 310.235 1286.070 310.605 ;
        RECT 1284.940 262.470 1285.080 310.235 ;
        RECT 1284.880 262.150 1285.140 262.470 ;
        RECT 1286.260 262.150 1286.520 262.470 ;
        RECT 1286.320 241.730 1286.460 262.150 ;
        RECT 1285.800 241.410 1286.060 241.730 ;
        RECT 1286.260 241.410 1286.520 241.730 ;
        RECT 1285.860 196.850 1286.000 241.410 ;
        RECT 1285.800 196.530 1286.060 196.850 ;
        RECT 1286.260 172.390 1286.520 172.710 ;
        RECT 1286.320 138.030 1286.460 172.390 ;
        RECT 1286.260 137.710 1286.520 138.030 ;
        RECT 1286.260 89.770 1286.520 90.090 ;
        RECT 1286.320 48.610 1286.460 89.770 ;
        RECT 1285.800 48.290 1286.060 48.610 ;
        RECT 1286.260 48.290 1286.520 48.610 ;
        RECT 1285.860 19.710 1286.000 48.290 ;
        RECT 1285.800 19.390 1286.060 19.710 ;
        RECT 1311.100 19.390 1311.360 19.710 ;
        RECT 1311.160 2.400 1311.300 19.390 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
      LAYER via2 ;
        RECT 1284.870 1296.960 1285.150 1297.240 ;
        RECT 1285.790 1296.960 1286.070 1297.240 ;
        RECT 1286.250 1145.320 1286.530 1145.600 ;
        RECT 1286.250 1144.640 1286.530 1144.920 ;
        RECT 1286.250 820.960 1286.530 821.240 ;
        RECT 1287.170 820.960 1287.450 821.240 ;
        RECT 1284.870 310.280 1285.150 310.560 ;
        RECT 1285.790 310.280 1286.070 310.560 ;
      LAYER met3 ;
        RECT 1284.845 1297.250 1285.175 1297.265 ;
        RECT 1285.765 1297.250 1286.095 1297.265 ;
        RECT 1284.845 1296.950 1286.095 1297.250 ;
        RECT 1284.845 1296.935 1285.175 1296.950 ;
        RECT 1285.765 1296.935 1286.095 1296.950 ;
        RECT 1286.225 1145.610 1286.555 1145.625 ;
        RECT 1285.550 1145.310 1286.555 1145.610 ;
        RECT 1285.550 1144.930 1285.850 1145.310 ;
        RECT 1286.225 1145.295 1286.555 1145.310 ;
        RECT 1286.225 1144.930 1286.555 1144.945 ;
        RECT 1285.550 1144.630 1286.555 1144.930 ;
        RECT 1286.225 1144.615 1286.555 1144.630 ;
        RECT 1286.225 821.250 1286.555 821.265 ;
        RECT 1287.145 821.250 1287.475 821.265 ;
        RECT 1286.225 820.950 1287.475 821.250 ;
        RECT 1286.225 820.935 1286.555 820.950 ;
        RECT 1287.145 820.935 1287.475 820.950 ;
        RECT 1284.845 310.570 1285.175 310.585 ;
        RECT 1285.765 310.570 1286.095 310.585 ;
        RECT 1284.845 310.270 1286.095 310.570 ;
        RECT 1284.845 310.255 1285.175 310.270 ;
        RECT 1285.765 310.255 1286.095 310.270 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1325.865 1676.625 1326.035 1687.335 ;
      LAYER mcon ;
        RECT 1325.865 1687.165 1326.035 1687.335 ;
      LAYER met1 ;
        RECT 1286.230 1687.320 1286.550 1687.380 ;
        RECT 1325.805 1687.320 1326.095 1687.365 ;
        RECT 1286.230 1687.180 1326.095 1687.320 ;
        RECT 1286.230 1687.120 1286.550 1687.180 ;
        RECT 1325.805 1687.135 1326.095 1687.180 ;
        RECT 1325.790 1676.780 1326.110 1676.840 ;
        RECT 1325.595 1676.640 1326.110 1676.780 ;
        RECT 1325.790 1676.580 1326.110 1676.640 ;
        RECT 1325.790 1635.300 1326.110 1635.360 ;
        RECT 1326.250 1635.300 1326.570 1635.360 ;
        RECT 1325.790 1635.160 1326.570 1635.300 ;
        RECT 1325.790 1635.100 1326.110 1635.160 ;
        RECT 1326.250 1635.100 1326.570 1635.160 ;
        RECT 1326.710 20.980 1327.030 21.040 ;
        RECT 1329.010 20.980 1329.330 21.040 ;
        RECT 1326.710 20.840 1329.330 20.980 ;
        RECT 1326.710 20.780 1327.030 20.840 ;
        RECT 1329.010 20.780 1329.330 20.840 ;
      LAYER via ;
        RECT 1286.260 1687.120 1286.520 1687.380 ;
        RECT 1325.820 1676.580 1326.080 1676.840 ;
        RECT 1325.820 1635.100 1326.080 1635.360 ;
        RECT 1326.280 1635.100 1326.540 1635.360 ;
        RECT 1326.740 20.780 1327.000 21.040 ;
        RECT 1329.040 20.780 1329.300 21.040 ;
      LAYER met2 ;
        RECT 1286.160 1700.340 1286.440 1704.000 ;
        RECT 1286.160 1700.000 1286.460 1700.340 ;
        RECT 1286.320 1687.410 1286.460 1700.000 ;
        RECT 1286.260 1687.090 1286.520 1687.410 ;
        RECT 1325.820 1676.550 1326.080 1676.870 ;
        RECT 1325.880 1635.390 1326.020 1676.550 ;
        RECT 1325.820 1635.070 1326.080 1635.390 ;
        RECT 1326.280 1635.070 1326.540 1635.390 ;
        RECT 1326.340 1514.770 1326.480 1635.070 ;
        RECT 1326.340 1514.630 1326.940 1514.770 ;
        RECT 1326.800 21.070 1326.940 1514.630 ;
        RECT 1326.740 20.750 1327.000 21.070 ;
        RECT 1329.040 20.750 1329.300 21.070 ;
        RECT 1329.100 2.400 1329.240 20.750 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 686.390 26.420 686.710 26.480 ;
        RECT 686.390 26.280 719.740 26.420 ;
        RECT 686.390 26.220 686.710 26.280 ;
        RECT 719.600 26.080 719.740 26.280 ;
        RECT 1219.990 26.080 1220.310 26.140 ;
        RECT 719.600 25.940 1220.310 26.080 ;
        RECT 1219.990 25.880 1220.310 25.940 ;
      LAYER via ;
        RECT 686.420 26.220 686.680 26.480 ;
        RECT 1220.020 25.880 1220.280 26.140 ;
      LAYER met2 ;
        RECT 1220.380 1700.410 1220.660 1704.000 ;
        RECT 1220.080 1700.270 1220.660 1700.410 ;
        RECT 686.420 26.190 686.680 26.510 ;
        RECT 686.480 2.400 686.620 26.190 ;
        RECT 1220.080 26.170 1220.220 1700.270 ;
        RECT 1220.380 1700.000 1220.660 1700.270 ;
        RECT 1220.020 25.850 1220.280 26.170 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1288.070 23.700 1288.390 23.760 ;
        RECT 1346.490 23.700 1346.810 23.760 ;
        RECT 1288.070 23.560 1346.810 23.700 ;
        RECT 1288.070 23.500 1288.390 23.560 ;
        RECT 1346.490 23.500 1346.810 23.560 ;
      LAYER via ;
        RECT 1288.100 23.500 1288.360 23.760 ;
        RECT 1346.520 23.500 1346.780 23.760 ;
      LAYER met2 ;
        RECT 1288.000 1700.340 1288.280 1704.000 ;
        RECT 1288.000 1700.000 1288.300 1700.340 ;
        RECT 1288.160 23.790 1288.300 1700.000 ;
        RECT 1288.100 23.470 1288.360 23.790 ;
        RECT 1346.520 23.470 1346.780 23.790 ;
        RECT 1346.580 2.400 1346.720 23.470 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1289.910 26.760 1290.230 26.820 ;
        RECT 1364.430 26.760 1364.750 26.820 ;
        RECT 1289.910 26.620 1364.750 26.760 ;
        RECT 1289.910 26.560 1290.230 26.620 ;
        RECT 1364.430 26.560 1364.750 26.620 ;
      LAYER via ;
        RECT 1289.940 26.560 1290.200 26.820 ;
        RECT 1364.460 26.560 1364.720 26.820 ;
      LAYER met2 ;
        RECT 1289.840 1700.340 1290.120 1704.000 ;
        RECT 1289.840 1700.000 1290.140 1700.340 ;
        RECT 1290.000 26.850 1290.140 1700.000 ;
        RECT 1289.940 26.530 1290.200 26.850 ;
        RECT 1364.460 26.530 1364.720 26.850 ;
        RECT 1364.520 2.400 1364.660 26.530 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1291.750 1678.820 1292.070 1678.880 ;
        RECT 1294.510 1678.820 1294.830 1678.880 ;
        RECT 1291.750 1678.680 1294.830 1678.820 ;
        RECT 1291.750 1678.620 1292.070 1678.680 ;
        RECT 1294.510 1678.620 1294.830 1678.680 ;
        RECT 1294.510 26.420 1294.830 26.480 ;
        RECT 1382.370 26.420 1382.690 26.480 ;
        RECT 1294.510 26.280 1382.690 26.420 ;
        RECT 1294.510 26.220 1294.830 26.280 ;
        RECT 1382.370 26.220 1382.690 26.280 ;
      LAYER via ;
        RECT 1291.780 1678.620 1292.040 1678.880 ;
        RECT 1294.540 1678.620 1294.800 1678.880 ;
        RECT 1294.540 26.220 1294.800 26.480 ;
        RECT 1382.400 26.220 1382.660 26.480 ;
      LAYER met2 ;
        RECT 1291.680 1700.340 1291.960 1704.000 ;
        RECT 1291.680 1700.000 1291.980 1700.340 ;
        RECT 1291.840 1678.910 1291.980 1700.000 ;
        RECT 1291.780 1678.590 1292.040 1678.910 ;
        RECT 1294.540 1678.590 1294.800 1678.910 ;
        RECT 1294.600 26.510 1294.740 1678.590 ;
        RECT 1294.540 26.190 1294.800 26.510 ;
        RECT 1382.400 26.190 1382.660 26.510 ;
        RECT 1382.460 2.400 1382.600 26.190 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1293.590 1683.920 1293.910 1683.980 ;
        RECT 1295.430 1683.920 1295.750 1683.980 ;
        RECT 1293.590 1683.780 1295.750 1683.920 ;
        RECT 1293.590 1683.720 1293.910 1683.780 ;
        RECT 1295.430 1683.720 1295.750 1683.780 ;
        RECT 1295.430 25.740 1295.750 25.800 ;
        RECT 1400.310 25.740 1400.630 25.800 ;
        RECT 1295.430 25.600 1400.630 25.740 ;
        RECT 1295.430 25.540 1295.750 25.600 ;
        RECT 1400.310 25.540 1400.630 25.600 ;
      LAYER via ;
        RECT 1293.620 1683.720 1293.880 1683.980 ;
        RECT 1295.460 1683.720 1295.720 1683.980 ;
        RECT 1295.460 25.540 1295.720 25.800 ;
        RECT 1400.340 25.540 1400.600 25.800 ;
      LAYER met2 ;
        RECT 1293.520 1700.340 1293.800 1704.000 ;
        RECT 1293.520 1700.000 1293.820 1700.340 ;
        RECT 1293.680 1684.010 1293.820 1700.000 ;
        RECT 1293.620 1683.690 1293.880 1684.010 ;
        RECT 1295.460 1683.690 1295.720 1684.010 ;
        RECT 1295.520 25.830 1295.660 1683.690 ;
        RECT 1295.460 25.510 1295.720 25.830 ;
        RECT 1400.340 25.510 1400.600 25.830 ;
        RECT 1400.400 2.400 1400.540 25.510 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1291.290 1684.600 1291.610 1684.660 ;
        RECT 1295.430 1684.600 1295.750 1684.660 ;
        RECT 1291.290 1684.460 1295.750 1684.600 ;
        RECT 1291.290 1684.400 1291.610 1684.460 ;
        RECT 1295.430 1684.400 1295.750 1684.460 ;
        RECT 1291.750 24.380 1292.070 24.440 ;
        RECT 1418.250 24.380 1418.570 24.440 ;
        RECT 1291.750 24.240 1418.570 24.380 ;
        RECT 1291.750 24.180 1292.070 24.240 ;
        RECT 1418.250 24.180 1418.570 24.240 ;
      LAYER via ;
        RECT 1291.320 1684.400 1291.580 1684.660 ;
        RECT 1295.460 1684.400 1295.720 1684.660 ;
        RECT 1291.780 24.180 1292.040 24.440 ;
        RECT 1418.280 24.180 1418.540 24.440 ;
      LAYER met2 ;
        RECT 1295.360 1700.340 1295.640 1704.000 ;
        RECT 1295.360 1700.000 1295.660 1700.340 ;
        RECT 1295.520 1684.690 1295.660 1700.000 ;
        RECT 1291.320 1684.370 1291.580 1684.690 ;
        RECT 1295.460 1684.370 1295.720 1684.690 ;
        RECT 1291.380 1678.140 1291.520 1684.370 ;
        RECT 1291.380 1678.000 1291.980 1678.140 ;
        RECT 1291.840 24.470 1291.980 1678.000 ;
        RECT 1291.780 24.150 1292.040 24.470 ;
        RECT 1418.280 24.150 1418.540 24.470 ;
        RECT 1418.340 2.400 1418.480 24.150 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1390.265 23.545 1390.435 24.735 ;
      LAYER mcon ;
        RECT 1390.265 24.565 1390.435 24.735 ;
      LAYER met1 ;
        RECT 1297.270 1683.920 1297.590 1683.980 ;
        RECT 1301.870 1683.920 1302.190 1683.980 ;
        RECT 1297.270 1683.780 1302.190 1683.920 ;
        RECT 1297.270 1683.720 1297.590 1683.780 ;
        RECT 1301.870 1683.720 1302.190 1683.780 ;
        RECT 1301.410 24.720 1301.730 24.780 ;
        RECT 1390.205 24.720 1390.495 24.765 ;
        RECT 1301.410 24.580 1390.495 24.720 ;
        RECT 1301.410 24.520 1301.730 24.580 ;
        RECT 1390.205 24.535 1390.495 24.580 ;
        RECT 1390.205 23.700 1390.495 23.745 ;
        RECT 1435.730 23.700 1436.050 23.760 ;
        RECT 1390.205 23.560 1436.050 23.700 ;
        RECT 1390.205 23.515 1390.495 23.560 ;
        RECT 1435.730 23.500 1436.050 23.560 ;
      LAYER via ;
        RECT 1297.300 1683.720 1297.560 1683.980 ;
        RECT 1301.900 1683.720 1302.160 1683.980 ;
        RECT 1301.440 24.520 1301.700 24.780 ;
        RECT 1435.760 23.500 1436.020 23.760 ;
      LAYER met2 ;
        RECT 1297.200 1700.340 1297.480 1704.000 ;
        RECT 1297.200 1700.000 1297.500 1700.340 ;
        RECT 1297.360 1684.010 1297.500 1700.000 ;
        RECT 1297.300 1683.690 1297.560 1684.010 ;
        RECT 1301.900 1683.690 1302.160 1684.010 ;
        RECT 1301.960 1677.290 1302.100 1683.690 ;
        RECT 1301.500 1677.150 1302.100 1677.290 ;
        RECT 1301.500 24.810 1301.640 1677.150 ;
        RECT 1301.440 24.490 1301.700 24.810 ;
        RECT 1435.760 23.470 1436.020 23.790 ;
        RECT 1435.820 2.400 1435.960 23.470 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1299.110 1666.920 1299.430 1666.980 ;
        RECT 1300.950 1666.920 1301.270 1666.980 ;
        RECT 1299.110 1666.780 1301.270 1666.920 ;
        RECT 1299.110 1666.720 1299.430 1666.780 ;
        RECT 1300.950 1666.720 1301.270 1666.780 ;
        RECT 1300.950 24.040 1301.270 24.100 ;
        RECT 1453.670 24.040 1453.990 24.100 ;
        RECT 1300.950 23.900 1453.990 24.040 ;
        RECT 1300.950 23.840 1301.270 23.900 ;
        RECT 1453.670 23.840 1453.990 23.900 ;
      LAYER via ;
        RECT 1299.140 1666.720 1299.400 1666.980 ;
        RECT 1300.980 1666.720 1301.240 1666.980 ;
        RECT 1300.980 23.840 1301.240 24.100 ;
        RECT 1453.700 23.840 1453.960 24.100 ;
      LAYER met2 ;
        RECT 1299.040 1700.340 1299.320 1704.000 ;
        RECT 1299.040 1700.000 1299.340 1700.340 ;
        RECT 1299.200 1667.010 1299.340 1700.000 ;
        RECT 1299.140 1666.690 1299.400 1667.010 ;
        RECT 1300.980 1666.690 1301.240 1667.010 ;
        RECT 1301.040 24.130 1301.180 1666.690 ;
        RECT 1300.980 23.810 1301.240 24.130 ;
        RECT 1453.700 23.810 1453.960 24.130 ;
        RECT 1453.760 2.400 1453.900 23.810 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1341.505 1685.125 1341.675 1688.015 ;
      LAYER mcon ;
        RECT 1341.505 1687.845 1341.675 1688.015 ;
      LAYER met1 ;
        RECT 1341.445 1688.000 1341.735 1688.045 ;
        RECT 1401.690 1688.000 1402.010 1688.060 ;
        RECT 1341.445 1687.860 1402.010 1688.000 ;
        RECT 1341.445 1687.815 1341.735 1687.860 ;
        RECT 1401.690 1687.800 1402.010 1687.860 ;
        RECT 1300.950 1685.280 1301.270 1685.340 ;
        RECT 1341.445 1685.280 1341.735 1685.325 ;
        RECT 1300.950 1685.140 1341.735 1685.280 ;
        RECT 1300.950 1685.080 1301.270 1685.140 ;
        RECT 1341.445 1685.095 1341.735 1685.140 ;
        RECT 1401.690 1683.240 1402.010 1683.300 ;
        RECT 1469.770 1683.240 1470.090 1683.300 ;
        RECT 1401.690 1683.100 1470.090 1683.240 ;
        RECT 1401.690 1683.040 1402.010 1683.100 ;
        RECT 1469.770 1683.040 1470.090 1683.100 ;
      LAYER via ;
        RECT 1401.720 1687.800 1401.980 1688.060 ;
        RECT 1300.980 1685.080 1301.240 1685.340 ;
        RECT 1401.720 1683.040 1401.980 1683.300 ;
        RECT 1469.800 1683.040 1470.060 1683.300 ;
      LAYER met2 ;
        RECT 1300.880 1700.340 1301.160 1704.000 ;
        RECT 1300.880 1700.000 1301.180 1700.340 ;
        RECT 1301.040 1685.370 1301.180 1700.000 ;
        RECT 1401.720 1687.770 1401.980 1688.090 ;
        RECT 1300.980 1685.050 1301.240 1685.370 ;
        RECT 1401.780 1683.330 1401.920 1687.770 ;
        RECT 1401.720 1683.010 1401.980 1683.330 ;
        RECT 1469.800 1683.010 1470.060 1683.330 ;
        RECT 1469.860 17.410 1470.000 1683.010 ;
        RECT 1469.860 17.270 1471.840 17.410 ;
        RECT 1471.700 2.400 1471.840 17.270 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1373.705 1682.745 1373.875 1687.675 ;
      LAYER mcon ;
        RECT 1373.705 1687.505 1373.875 1687.675 ;
      LAYER met1 ;
        RECT 1327.720 1687.860 1337.980 1688.000 ;
        RECT 1302.790 1686.980 1303.110 1687.040 ;
        RECT 1327.720 1686.980 1327.860 1687.860 ;
        RECT 1337.840 1687.660 1337.980 1687.860 ;
        RECT 1373.645 1687.660 1373.935 1687.705 ;
        RECT 1337.840 1687.520 1373.935 1687.660 ;
        RECT 1373.645 1687.475 1373.935 1687.520 ;
        RECT 1302.790 1686.840 1327.860 1686.980 ;
        RECT 1302.790 1686.780 1303.110 1686.840 ;
        RECT 1373.645 1682.900 1373.935 1682.945 ;
        RECT 1483.570 1682.900 1483.890 1682.960 ;
        RECT 1373.645 1682.760 1483.890 1682.900 ;
        RECT 1373.645 1682.715 1373.935 1682.760 ;
        RECT 1483.570 1682.700 1483.890 1682.760 ;
        RECT 1483.570 20.980 1483.890 21.040 ;
        RECT 1489.550 20.980 1489.870 21.040 ;
        RECT 1483.570 20.840 1489.870 20.980 ;
        RECT 1483.570 20.780 1483.890 20.840 ;
        RECT 1489.550 20.780 1489.870 20.840 ;
      LAYER via ;
        RECT 1302.820 1686.780 1303.080 1687.040 ;
        RECT 1483.600 1682.700 1483.860 1682.960 ;
        RECT 1483.600 20.780 1483.860 21.040 ;
        RECT 1489.580 20.780 1489.840 21.040 ;
      LAYER met2 ;
        RECT 1302.720 1700.340 1303.000 1704.000 ;
        RECT 1302.720 1700.000 1303.020 1700.340 ;
        RECT 1302.880 1687.070 1303.020 1700.000 ;
        RECT 1302.820 1686.750 1303.080 1687.070 ;
        RECT 1483.600 1682.670 1483.860 1682.990 ;
        RECT 1483.660 21.070 1483.800 1682.670 ;
        RECT 1483.600 20.750 1483.860 21.070 ;
        RECT 1489.580 20.750 1489.840 21.070 ;
        RECT 1489.640 2.400 1489.780 20.750 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1449.145 1679.685 1449.315 1682.575 ;
      LAYER mcon ;
        RECT 1449.145 1682.405 1449.315 1682.575 ;
      LAYER met1 ;
        RECT 1304.630 1682.560 1304.950 1682.620 ;
        RECT 1449.085 1682.560 1449.375 1682.605 ;
        RECT 1304.630 1682.420 1449.375 1682.560 ;
        RECT 1304.630 1682.360 1304.950 1682.420 ;
        RECT 1449.085 1682.375 1449.375 1682.420 ;
        RECT 1449.085 1679.840 1449.375 1679.885 ;
        RECT 1504.270 1679.840 1504.590 1679.900 ;
        RECT 1449.085 1679.700 1504.590 1679.840 ;
        RECT 1449.085 1679.655 1449.375 1679.700 ;
        RECT 1504.270 1679.640 1504.590 1679.700 ;
        RECT 1504.270 2.960 1504.590 3.020 ;
        RECT 1507.030 2.960 1507.350 3.020 ;
        RECT 1504.270 2.820 1507.350 2.960 ;
        RECT 1504.270 2.760 1504.590 2.820 ;
        RECT 1507.030 2.760 1507.350 2.820 ;
      LAYER via ;
        RECT 1304.660 1682.360 1304.920 1682.620 ;
        RECT 1504.300 1679.640 1504.560 1679.900 ;
        RECT 1504.300 2.760 1504.560 3.020 ;
        RECT 1507.060 2.760 1507.320 3.020 ;
      LAYER met2 ;
        RECT 1304.560 1700.340 1304.840 1704.000 ;
        RECT 1304.560 1700.000 1304.860 1700.340 ;
        RECT 1304.720 1682.650 1304.860 1700.000 ;
        RECT 1304.660 1682.330 1304.920 1682.650 ;
        RECT 1504.300 1679.610 1504.560 1679.930 ;
        RECT 1504.360 3.050 1504.500 1679.610 ;
        RECT 1504.300 2.730 1504.560 3.050 ;
        RECT 1507.060 2.730 1507.320 3.050 ;
        RECT 1507.120 2.400 1507.260 2.730 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 710.310 1667.260 710.630 1667.320 ;
        RECT 1222.290 1667.260 1222.610 1667.320 ;
        RECT 710.310 1667.120 1222.610 1667.260 ;
        RECT 710.310 1667.060 710.630 1667.120 ;
        RECT 1222.290 1667.060 1222.610 1667.120 ;
        RECT 704.330 26.080 704.650 26.140 ;
        RECT 710.310 26.080 710.630 26.140 ;
        RECT 704.330 25.940 710.630 26.080 ;
        RECT 704.330 25.880 704.650 25.940 ;
        RECT 710.310 25.880 710.630 25.940 ;
      LAYER via ;
        RECT 710.340 1667.060 710.600 1667.320 ;
        RECT 1222.320 1667.060 1222.580 1667.320 ;
        RECT 704.360 25.880 704.620 26.140 ;
        RECT 710.340 25.880 710.600 26.140 ;
      LAYER met2 ;
        RECT 1222.220 1700.340 1222.500 1704.000 ;
        RECT 1222.220 1700.000 1222.520 1700.340 ;
        RECT 1222.380 1667.350 1222.520 1700.000 ;
        RECT 710.340 1667.030 710.600 1667.350 ;
        RECT 1222.320 1667.030 1222.580 1667.350 ;
        RECT 710.400 26.170 710.540 1667.030 ;
        RECT 704.360 25.850 704.620 26.170 ;
        RECT 710.340 25.850 710.600 26.170 ;
        RECT 704.420 2.400 704.560 25.850 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1341.965 1689.205 1342.135 1690.395 ;
        RECT 1389.345 1686.485 1389.515 1688.695 ;
      LAYER mcon ;
        RECT 1341.965 1690.225 1342.135 1690.395 ;
        RECT 1389.345 1688.525 1389.515 1688.695 ;
      LAYER met1 ;
        RECT 1306.470 1690.380 1306.790 1690.440 ;
        RECT 1341.905 1690.380 1342.195 1690.425 ;
        RECT 1306.470 1690.240 1342.195 1690.380 ;
        RECT 1306.470 1690.180 1306.790 1690.240 ;
        RECT 1341.905 1690.195 1342.195 1690.240 ;
        RECT 1341.905 1689.360 1342.195 1689.405 ;
        RECT 1341.905 1689.220 1363.740 1689.360 ;
        RECT 1341.905 1689.175 1342.195 1689.220 ;
        RECT 1363.600 1688.680 1363.740 1689.220 ;
        RECT 1389.285 1688.680 1389.575 1688.725 ;
        RECT 1363.600 1688.540 1389.575 1688.680 ;
        RECT 1389.285 1688.495 1389.575 1688.540 ;
        RECT 1389.285 1686.640 1389.575 1686.685 ;
        RECT 1405.370 1686.640 1405.690 1686.700 ;
        RECT 1389.285 1686.500 1405.690 1686.640 ;
        RECT 1389.285 1686.455 1389.575 1686.500 ;
        RECT 1405.370 1686.440 1405.690 1686.500 ;
        RECT 1405.370 1675.760 1405.690 1675.820 ;
        RECT 1524.970 1675.760 1525.290 1675.820 ;
        RECT 1405.370 1675.620 1525.290 1675.760 ;
        RECT 1405.370 1675.560 1405.690 1675.620 ;
        RECT 1524.970 1675.560 1525.290 1675.620 ;
      LAYER via ;
        RECT 1306.500 1690.180 1306.760 1690.440 ;
        RECT 1405.400 1686.440 1405.660 1686.700 ;
        RECT 1405.400 1675.560 1405.660 1675.820 ;
        RECT 1525.000 1675.560 1525.260 1675.820 ;
      LAYER met2 ;
        RECT 1306.400 1700.340 1306.680 1704.000 ;
        RECT 1306.400 1700.000 1306.700 1700.340 ;
        RECT 1306.560 1690.470 1306.700 1700.000 ;
        RECT 1306.500 1690.150 1306.760 1690.470 ;
        RECT 1405.400 1686.410 1405.660 1686.730 ;
        RECT 1405.460 1675.850 1405.600 1686.410 ;
        RECT 1405.400 1675.530 1405.660 1675.850 ;
        RECT 1525.000 1675.530 1525.260 1675.850 ;
        RECT 1525.060 2.400 1525.200 1675.530 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1393.945 1668.465 1394.115 1669.995 ;
        RECT 1441.785 1668.805 1441.955 1669.995 ;
        RECT 1490.545 1668.465 1490.715 1669.995 ;
        RECT 1538.385 1669.145 1538.555 1669.995 ;
      LAYER mcon ;
        RECT 1393.945 1669.825 1394.115 1669.995 ;
        RECT 1441.785 1669.825 1441.955 1669.995 ;
        RECT 1490.545 1669.825 1490.715 1669.995 ;
        RECT 1538.385 1669.825 1538.555 1669.995 ;
      LAYER met1 ;
        RECT 1393.885 1669.980 1394.175 1670.025 ;
        RECT 1441.725 1669.980 1442.015 1670.025 ;
        RECT 1393.885 1669.840 1442.015 1669.980 ;
        RECT 1393.885 1669.795 1394.175 1669.840 ;
        RECT 1441.725 1669.795 1442.015 1669.840 ;
        RECT 1490.485 1669.980 1490.775 1670.025 ;
        RECT 1538.325 1669.980 1538.615 1670.025 ;
        RECT 1490.485 1669.840 1538.615 1669.980 ;
        RECT 1490.485 1669.795 1490.775 1669.840 ;
        RECT 1538.325 1669.795 1538.615 1669.840 ;
        RECT 1538.325 1669.115 1538.615 1669.345 ;
        RECT 1308.310 1668.760 1308.630 1669.020 ;
        RECT 1441.725 1668.775 1442.015 1669.005 ;
        RECT 1538.400 1668.960 1538.540 1669.115 ;
        RECT 1538.770 1668.960 1539.090 1669.020 ;
        RECT 1538.400 1668.820 1539.090 1668.960 ;
        RECT 1308.400 1668.620 1308.540 1668.760 ;
        RECT 1393.885 1668.620 1394.175 1668.665 ;
        RECT 1308.400 1668.480 1394.175 1668.620 ;
        RECT 1441.800 1668.620 1441.940 1668.775 ;
        RECT 1538.770 1668.760 1539.090 1668.820 ;
        RECT 1490.485 1668.620 1490.775 1668.665 ;
        RECT 1441.800 1668.480 1490.775 1668.620 ;
        RECT 1393.885 1668.435 1394.175 1668.480 ;
        RECT 1490.485 1668.435 1490.775 1668.480 ;
      LAYER via ;
        RECT 1308.340 1668.760 1308.600 1669.020 ;
        RECT 1538.800 1668.760 1539.060 1669.020 ;
      LAYER met2 ;
        RECT 1308.240 1700.340 1308.520 1704.000 ;
        RECT 1308.240 1700.000 1308.540 1700.340 ;
        RECT 1308.400 1669.050 1308.540 1700.000 ;
        RECT 1308.340 1668.730 1308.600 1669.050 ;
        RECT 1538.790 1668.705 1539.070 1669.075 ;
        RECT 1538.790 1667.515 1539.070 1667.885 ;
        RECT 1538.860 17.410 1539.000 1667.515 ;
        RECT 1538.860 17.270 1543.140 17.410 ;
        RECT 1543.000 2.400 1543.140 17.270 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
      LAYER via2 ;
        RECT 1538.790 1668.750 1539.070 1669.030 ;
        RECT 1538.790 1667.560 1539.070 1667.840 ;
      LAYER met3 ;
        RECT 1538.765 1669.040 1539.095 1669.055 ;
        RECT 1538.550 1668.725 1539.095 1669.040 ;
        RECT 1538.550 1667.865 1538.850 1668.725 ;
        RECT 1538.550 1667.550 1539.095 1667.865 ;
        RECT 1538.765 1667.535 1539.095 1667.550 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1310.150 1675.080 1310.470 1675.140 ;
        RECT 1559.470 1675.080 1559.790 1675.140 ;
        RECT 1310.150 1674.940 1559.790 1675.080 ;
        RECT 1310.150 1674.880 1310.470 1674.940 ;
        RECT 1559.470 1674.880 1559.790 1674.940 ;
      LAYER via ;
        RECT 1310.180 1674.880 1310.440 1675.140 ;
        RECT 1559.500 1674.880 1559.760 1675.140 ;
      LAYER met2 ;
        RECT 1310.080 1700.340 1310.360 1704.000 ;
        RECT 1310.080 1700.000 1310.380 1700.340 ;
        RECT 1310.240 1675.170 1310.380 1700.000 ;
        RECT 1310.180 1674.850 1310.440 1675.170 ;
        RECT 1559.500 1674.850 1559.760 1675.170 ;
        RECT 1559.560 17.410 1559.700 1674.850 ;
        RECT 1559.560 17.270 1561.080 17.410 ;
        RECT 1560.940 2.400 1561.080 17.270 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1312.450 1682.220 1312.770 1682.280 ;
        RECT 1573.270 1682.220 1573.590 1682.280 ;
        RECT 1312.450 1682.080 1573.590 1682.220 ;
        RECT 1312.450 1682.020 1312.770 1682.080 ;
        RECT 1573.270 1682.020 1573.590 1682.080 ;
      LAYER via ;
        RECT 1312.480 1682.020 1312.740 1682.280 ;
        RECT 1573.300 1682.020 1573.560 1682.280 ;
      LAYER met2 ;
        RECT 1311.920 1700.340 1312.200 1704.000 ;
        RECT 1311.920 1700.000 1312.220 1700.340 ;
        RECT 1312.080 1685.450 1312.220 1700.000 ;
        RECT 1312.080 1685.310 1312.680 1685.450 ;
        RECT 1312.540 1682.310 1312.680 1685.310 ;
        RECT 1312.480 1681.990 1312.740 1682.310 ;
        RECT 1573.300 1681.990 1573.560 1682.310 ;
        RECT 1573.360 18.090 1573.500 1681.990 ;
        RECT 1573.360 17.950 1579.020 18.090 ;
        RECT 1578.880 2.400 1579.020 17.950 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1376.465 1689.205 1376.635 1690.055 ;
      LAYER mcon ;
        RECT 1376.465 1689.885 1376.635 1690.055 ;
      LAYER met1 ;
        RECT 1313.830 1690.040 1314.150 1690.100 ;
        RECT 1376.405 1690.040 1376.695 1690.085 ;
        RECT 1403.530 1690.040 1403.850 1690.100 ;
        RECT 1313.830 1689.900 1365.120 1690.040 ;
        RECT 1313.830 1689.840 1314.150 1689.900 ;
        RECT 1364.980 1689.360 1365.120 1689.900 ;
        RECT 1376.405 1689.900 1403.850 1690.040 ;
        RECT 1376.405 1689.855 1376.695 1689.900 ;
        RECT 1403.530 1689.840 1403.850 1689.900 ;
        RECT 1376.405 1689.360 1376.695 1689.405 ;
        RECT 1364.980 1689.220 1376.695 1689.360 ;
        RECT 1376.405 1689.175 1376.695 1689.220 ;
        RECT 1403.530 1685.960 1403.850 1686.020 ;
        RECT 1405.830 1685.960 1406.150 1686.020 ;
        RECT 1403.530 1685.820 1406.150 1685.960 ;
        RECT 1403.530 1685.760 1403.850 1685.820 ;
        RECT 1405.830 1685.760 1406.150 1685.820 ;
        RECT 1405.830 1661.480 1406.150 1661.540 ;
        RECT 1593.970 1661.480 1594.290 1661.540 ;
        RECT 1405.830 1661.340 1594.290 1661.480 ;
        RECT 1405.830 1661.280 1406.150 1661.340 ;
        RECT 1593.970 1661.280 1594.290 1661.340 ;
      LAYER via ;
        RECT 1313.860 1689.840 1314.120 1690.100 ;
        RECT 1403.560 1689.840 1403.820 1690.100 ;
        RECT 1403.560 1685.760 1403.820 1686.020 ;
        RECT 1405.860 1685.760 1406.120 1686.020 ;
        RECT 1405.860 1661.280 1406.120 1661.540 ;
        RECT 1594.000 1661.280 1594.260 1661.540 ;
      LAYER met2 ;
        RECT 1313.760 1700.340 1314.040 1704.000 ;
        RECT 1313.760 1700.000 1314.060 1700.340 ;
        RECT 1313.920 1690.130 1314.060 1700.000 ;
        RECT 1313.860 1689.810 1314.120 1690.130 ;
        RECT 1403.560 1689.810 1403.820 1690.130 ;
        RECT 1403.620 1686.050 1403.760 1689.810 ;
        RECT 1403.560 1685.730 1403.820 1686.050 ;
        RECT 1405.860 1685.730 1406.120 1686.050 ;
        RECT 1405.920 1661.570 1406.060 1685.730 ;
        RECT 1405.860 1661.250 1406.120 1661.570 ;
        RECT 1594.000 1661.250 1594.260 1661.570 ;
        RECT 1594.060 17.410 1594.200 1661.250 ;
        RECT 1594.060 17.270 1596.500 17.410 ;
        RECT 1596.360 2.400 1596.500 17.270 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1313.830 1683.920 1314.150 1683.980 ;
        RECT 1315.670 1683.920 1315.990 1683.980 ;
        RECT 1313.830 1683.780 1315.990 1683.920 ;
        RECT 1313.830 1683.720 1314.150 1683.780 ;
        RECT 1315.670 1683.720 1315.990 1683.780 ;
        RECT 1313.830 27.780 1314.150 27.840 ;
        RECT 1614.210 27.780 1614.530 27.840 ;
        RECT 1313.830 27.640 1614.530 27.780 ;
        RECT 1313.830 27.580 1314.150 27.640 ;
        RECT 1614.210 27.580 1614.530 27.640 ;
      LAYER via ;
        RECT 1313.860 1683.720 1314.120 1683.980 ;
        RECT 1315.700 1683.720 1315.960 1683.980 ;
        RECT 1313.860 27.580 1314.120 27.840 ;
        RECT 1614.240 27.580 1614.500 27.840 ;
      LAYER met2 ;
        RECT 1315.600 1700.340 1315.880 1704.000 ;
        RECT 1315.600 1700.000 1315.900 1700.340 ;
        RECT 1315.760 1684.010 1315.900 1700.000 ;
        RECT 1313.860 1683.690 1314.120 1684.010 ;
        RECT 1315.700 1683.690 1315.960 1684.010 ;
        RECT 1313.920 27.870 1314.060 1683.690 ;
        RECT 1313.860 27.550 1314.120 27.870 ;
        RECT 1614.240 27.550 1614.500 27.870 ;
        RECT 1614.300 2.400 1614.440 27.550 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1312.525 1145.205 1312.695 1173.595 ;
        RECT 1313.445 993.565 1313.615 1089.955 ;
        RECT 1313.445 897.005 1313.615 945.115 ;
        RECT 1313.445 800.445 1313.615 848.555 ;
        RECT 1313.445 655.605 1313.615 703.715 ;
        RECT 1313.445 511.105 1313.615 558.875 ;
        RECT 1313.445 455.345 1313.615 510.595 ;
        RECT 1312.985 34.765 1313.155 82.875 ;
      LAYER mcon ;
        RECT 1312.525 1173.425 1312.695 1173.595 ;
        RECT 1313.445 1089.785 1313.615 1089.955 ;
        RECT 1313.445 944.945 1313.615 945.115 ;
        RECT 1313.445 848.385 1313.615 848.555 ;
        RECT 1313.445 703.545 1313.615 703.715 ;
        RECT 1313.445 558.705 1313.615 558.875 ;
        RECT 1313.445 510.425 1313.615 510.595 ;
        RECT 1312.985 82.705 1313.155 82.875 ;
      LAYER met1 ;
        RECT 1313.370 1621.700 1313.690 1621.760 ;
        RECT 1317.970 1621.700 1318.290 1621.760 ;
        RECT 1313.370 1621.560 1318.290 1621.700 ;
        RECT 1313.370 1621.500 1313.690 1621.560 ;
        RECT 1317.970 1621.500 1318.290 1621.560 ;
        RECT 1311.990 1573.420 1312.310 1573.480 ;
        RECT 1312.910 1573.420 1313.230 1573.480 ;
        RECT 1311.990 1573.280 1313.230 1573.420 ;
        RECT 1311.990 1573.220 1312.310 1573.280 ;
        RECT 1312.910 1573.220 1313.230 1573.280 ;
        RECT 1312.910 1532.620 1313.230 1532.680 ;
        RECT 1312.910 1532.480 1313.600 1532.620 ;
        RECT 1312.910 1532.420 1313.230 1532.480 ;
        RECT 1313.460 1532.000 1313.600 1532.480 ;
        RECT 1313.370 1531.740 1313.690 1532.000 ;
        RECT 1312.450 1235.120 1312.770 1235.180 ;
        RECT 1313.370 1235.120 1313.690 1235.180 ;
        RECT 1312.450 1234.980 1313.690 1235.120 ;
        RECT 1312.450 1234.920 1312.770 1234.980 ;
        RECT 1313.370 1234.920 1313.690 1234.980 ;
        RECT 1312.465 1173.580 1312.755 1173.625 ;
        RECT 1313.370 1173.580 1313.690 1173.640 ;
        RECT 1312.465 1173.440 1313.690 1173.580 ;
        RECT 1312.465 1173.395 1312.755 1173.440 ;
        RECT 1313.370 1173.380 1313.690 1173.440 ;
        RECT 1312.450 1145.360 1312.770 1145.420 ;
        RECT 1312.255 1145.220 1312.770 1145.360 ;
        RECT 1312.450 1145.160 1312.770 1145.220 ;
        RECT 1313.370 1089.940 1313.690 1090.000 ;
        RECT 1313.175 1089.800 1313.690 1089.940 ;
        RECT 1313.370 1089.740 1313.690 1089.800 ;
        RECT 1313.370 993.720 1313.690 993.780 ;
        RECT 1313.175 993.580 1313.690 993.720 ;
        RECT 1313.370 993.520 1313.690 993.580 ;
        RECT 1313.370 945.100 1313.690 945.160 ;
        RECT 1313.175 944.960 1313.690 945.100 ;
        RECT 1313.370 944.900 1313.690 944.960 ;
        RECT 1313.370 897.160 1313.690 897.220 ;
        RECT 1313.175 897.020 1313.690 897.160 ;
        RECT 1313.370 896.960 1313.690 897.020 ;
        RECT 1313.370 848.540 1313.690 848.600 ;
        RECT 1313.175 848.400 1313.690 848.540 ;
        RECT 1313.370 848.340 1313.690 848.400 ;
        RECT 1313.370 800.600 1313.690 800.660 ;
        RECT 1313.175 800.460 1313.690 800.600 ;
        RECT 1313.370 800.400 1313.690 800.460 ;
        RECT 1313.370 703.700 1313.690 703.760 ;
        RECT 1313.175 703.560 1313.690 703.700 ;
        RECT 1313.370 703.500 1313.690 703.560 ;
        RECT 1313.370 655.760 1313.690 655.820 ;
        RECT 1313.175 655.620 1313.690 655.760 ;
        RECT 1313.370 655.560 1313.690 655.620 ;
        RECT 1313.370 558.860 1313.690 558.920 ;
        RECT 1313.175 558.720 1313.690 558.860 ;
        RECT 1313.370 558.660 1313.690 558.720 ;
        RECT 1313.370 511.260 1313.690 511.320 ;
        RECT 1313.175 511.120 1313.690 511.260 ;
        RECT 1313.370 511.060 1313.690 511.120 ;
        RECT 1313.370 510.580 1313.690 510.640 ;
        RECT 1313.175 510.440 1313.690 510.580 ;
        RECT 1313.370 510.380 1313.690 510.440 ;
        RECT 1312.910 455.500 1313.230 455.560 ;
        RECT 1313.385 455.500 1313.675 455.545 ;
        RECT 1312.910 455.360 1313.675 455.500 ;
        RECT 1312.910 455.300 1313.230 455.360 ;
        RECT 1313.385 455.315 1313.675 455.360 ;
        RECT 1312.910 407.220 1313.230 407.280 ;
        RECT 1312.540 407.080 1313.230 407.220 ;
        RECT 1312.540 406.940 1312.680 407.080 ;
        RECT 1312.910 407.020 1313.230 407.080 ;
        RECT 1312.450 406.680 1312.770 406.940 ;
        RECT 1312.910 227.700 1313.230 227.760 ;
        RECT 1313.370 227.700 1313.690 227.760 ;
        RECT 1312.910 227.560 1313.690 227.700 ;
        RECT 1312.910 227.500 1313.230 227.560 ;
        RECT 1313.370 227.500 1313.690 227.560 ;
        RECT 1312.925 82.860 1313.215 82.905 ;
        RECT 1313.370 82.860 1313.690 82.920 ;
        RECT 1312.925 82.720 1313.690 82.860 ;
        RECT 1312.925 82.675 1313.215 82.720 ;
        RECT 1313.370 82.660 1313.690 82.720 ;
        RECT 1312.910 34.920 1313.230 34.980 ;
        RECT 1312.715 34.780 1313.230 34.920 ;
        RECT 1312.910 34.720 1313.230 34.780 ;
        RECT 1313.370 28.120 1313.690 28.180 ;
        RECT 1632.150 28.120 1632.470 28.180 ;
        RECT 1313.370 27.980 1632.470 28.120 ;
        RECT 1313.370 27.920 1313.690 27.980 ;
        RECT 1632.150 27.920 1632.470 27.980 ;
      LAYER via ;
        RECT 1313.400 1621.500 1313.660 1621.760 ;
        RECT 1318.000 1621.500 1318.260 1621.760 ;
        RECT 1312.020 1573.220 1312.280 1573.480 ;
        RECT 1312.940 1573.220 1313.200 1573.480 ;
        RECT 1312.940 1532.420 1313.200 1532.680 ;
        RECT 1313.400 1531.740 1313.660 1532.000 ;
        RECT 1312.480 1234.920 1312.740 1235.180 ;
        RECT 1313.400 1234.920 1313.660 1235.180 ;
        RECT 1313.400 1173.380 1313.660 1173.640 ;
        RECT 1312.480 1145.160 1312.740 1145.420 ;
        RECT 1313.400 1089.740 1313.660 1090.000 ;
        RECT 1313.400 993.520 1313.660 993.780 ;
        RECT 1313.400 944.900 1313.660 945.160 ;
        RECT 1313.400 896.960 1313.660 897.220 ;
        RECT 1313.400 848.340 1313.660 848.600 ;
        RECT 1313.400 800.400 1313.660 800.660 ;
        RECT 1313.400 703.500 1313.660 703.760 ;
        RECT 1313.400 655.560 1313.660 655.820 ;
        RECT 1313.400 558.660 1313.660 558.920 ;
        RECT 1313.400 511.060 1313.660 511.320 ;
        RECT 1313.400 510.380 1313.660 510.640 ;
        RECT 1312.940 455.300 1313.200 455.560 ;
        RECT 1312.940 407.020 1313.200 407.280 ;
        RECT 1312.480 406.680 1312.740 406.940 ;
        RECT 1312.940 227.500 1313.200 227.760 ;
        RECT 1313.400 227.500 1313.660 227.760 ;
        RECT 1313.400 82.660 1313.660 82.920 ;
        RECT 1312.940 34.720 1313.200 34.980 ;
        RECT 1313.400 27.920 1313.660 28.180 ;
        RECT 1632.180 27.920 1632.440 28.180 ;
      LAYER met2 ;
        RECT 1317.440 1700.340 1317.720 1704.000 ;
        RECT 1317.440 1700.000 1317.740 1700.340 ;
        RECT 1317.600 1691.570 1317.740 1700.000 ;
        RECT 1317.600 1691.430 1318.200 1691.570 ;
        RECT 1318.060 1621.790 1318.200 1691.430 ;
        RECT 1313.400 1621.645 1313.660 1621.790 ;
        RECT 1312.010 1621.275 1312.290 1621.645 ;
        RECT 1313.390 1621.275 1313.670 1621.645 ;
        RECT 1318.000 1621.470 1318.260 1621.790 ;
        RECT 1312.080 1573.510 1312.220 1621.275 ;
        RECT 1312.020 1573.190 1312.280 1573.510 ;
        RECT 1312.940 1573.190 1313.200 1573.510 ;
        RECT 1313.000 1532.710 1313.140 1573.190 ;
        RECT 1312.940 1532.390 1313.200 1532.710 ;
        RECT 1313.400 1531.710 1313.660 1532.030 ;
        RECT 1313.460 1332.530 1313.600 1531.710 ;
        RECT 1313.000 1332.390 1313.600 1332.530 ;
        RECT 1313.000 1331.850 1313.140 1332.390 ;
        RECT 1313.000 1331.710 1313.600 1331.850 ;
        RECT 1313.460 1235.210 1313.600 1331.710 ;
        RECT 1312.480 1234.890 1312.740 1235.210 ;
        RECT 1313.400 1234.890 1313.660 1235.210 ;
        RECT 1312.540 1187.125 1312.680 1234.890 ;
        RECT 1312.470 1186.755 1312.750 1187.125 ;
        RECT 1313.390 1186.755 1313.670 1187.125 ;
        RECT 1313.460 1173.670 1313.600 1186.755 ;
        RECT 1313.400 1173.350 1313.660 1173.670 ;
        RECT 1312.480 1145.130 1312.740 1145.450 ;
        RECT 1312.540 1097.250 1312.680 1145.130 ;
        RECT 1312.540 1097.110 1313.600 1097.250 ;
        RECT 1313.460 1090.030 1313.600 1097.110 ;
        RECT 1313.400 1089.710 1313.660 1090.030 ;
        RECT 1313.400 993.490 1313.660 993.810 ;
        RECT 1313.460 945.190 1313.600 993.490 ;
        RECT 1313.400 944.870 1313.660 945.190 ;
        RECT 1313.400 896.930 1313.660 897.250 ;
        RECT 1313.460 848.630 1313.600 896.930 ;
        RECT 1313.400 848.310 1313.660 848.630 ;
        RECT 1313.400 800.370 1313.660 800.690 ;
        RECT 1313.460 703.790 1313.600 800.370 ;
        RECT 1313.400 703.470 1313.660 703.790 ;
        RECT 1313.400 655.530 1313.660 655.850 ;
        RECT 1313.460 558.950 1313.600 655.530 ;
        RECT 1313.400 558.630 1313.660 558.950 ;
        RECT 1313.400 511.030 1313.660 511.350 ;
        RECT 1313.460 510.670 1313.600 511.030 ;
        RECT 1313.400 510.350 1313.660 510.670 ;
        RECT 1312.940 455.270 1313.200 455.590 ;
        RECT 1313.000 407.310 1313.140 455.270 ;
        RECT 1312.940 406.990 1313.200 407.310 ;
        RECT 1312.480 406.650 1312.740 406.970 ;
        RECT 1312.540 376.450 1312.680 406.650 ;
        RECT 1312.080 376.310 1312.680 376.450 ;
        RECT 1312.080 334.290 1312.220 376.310 ;
        RECT 1312.080 334.150 1313.140 334.290 ;
        RECT 1313.000 227.790 1313.140 334.150 ;
        RECT 1312.940 227.470 1313.200 227.790 ;
        RECT 1313.400 227.470 1313.660 227.790 ;
        RECT 1313.460 82.950 1313.600 227.470 ;
        RECT 1313.400 82.630 1313.660 82.950 ;
        RECT 1312.940 34.690 1313.200 35.010 ;
        RECT 1313.000 34.240 1313.140 34.690 ;
        RECT 1313.000 34.100 1313.600 34.240 ;
        RECT 1313.460 28.210 1313.600 34.100 ;
        RECT 1313.400 27.890 1313.660 28.210 ;
        RECT 1632.180 27.890 1632.440 28.210 ;
        RECT 1632.240 2.400 1632.380 27.890 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
      LAYER via2 ;
        RECT 1312.010 1621.320 1312.290 1621.600 ;
        RECT 1313.390 1621.320 1313.670 1621.600 ;
        RECT 1312.470 1186.800 1312.750 1187.080 ;
        RECT 1313.390 1186.800 1313.670 1187.080 ;
      LAYER met3 ;
        RECT 1311.985 1621.610 1312.315 1621.625 ;
        RECT 1313.365 1621.610 1313.695 1621.625 ;
        RECT 1311.985 1621.310 1313.695 1621.610 ;
        RECT 1311.985 1621.295 1312.315 1621.310 ;
        RECT 1313.365 1621.295 1313.695 1621.310 ;
        RECT 1312.445 1187.090 1312.775 1187.105 ;
        RECT 1313.365 1187.090 1313.695 1187.105 ;
        RECT 1312.445 1186.790 1313.695 1187.090 ;
        RECT 1312.445 1186.775 1312.775 1186.790 ;
        RECT 1313.365 1186.775 1313.695 1186.790 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1321.265 1097.265 1321.435 1186.855 ;
        RECT 1321.265 1041.845 1321.435 1089.955 ;
        RECT 1321.265 897.005 1321.435 945.115 ;
        RECT 1321.265 800.445 1321.435 848.555 ;
        RECT 1321.265 655.605 1321.435 703.715 ;
        RECT 1321.265 462.485 1321.435 510.595 ;
        RECT 1321.265 378.845 1321.435 414.035 ;
        RECT 1321.265 179.605 1321.435 227.715 ;
        RECT 1321.265 83.045 1321.435 131.155 ;
        RECT 1321.265 28.305 1321.435 34.255 ;
      LAYER mcon ;
        RECT 1321.265 1186.685 1321.435 1186.855 ;
        RECT 1321.265 1089.785 1321.435 1089.955 ;
        RECT 1321.265 944.945 1321.435 945.115 ;
        RECT 1321.265 848.385 1321.435 848.555 ;
        RECT 1321.265 703.545 1321.435 703.715 ;
        RECT 1321.265 510.425 1321.435 510.595 ;
        RECT 1321.265 413.865 1321.435 414.035 ;
        RECT 1321.265 227.545 1321.435 227.715 ;
        RECT 1321.265 130.985 1321.435 131.155 ;
        RECT 1321.265 34.085 1321.435 34.255 ;
      LAYER met1 ;
        RECT 1319.350 1634.960 1319.670 1635.020 ;
        RECT 1321.650 1634.960 1321.970 1635.020 ;
        RECT 1319.350 1634.820 1321.970 1634.960 ;
        RECT 1319.350 1634.760 1319.670 1634.820 ;
        RECT 1321.650 1634.760 1321.970 1634.820 ;
        RECT 1321.190 1531.940 1321.510 1532.000 ;
        RECT 1321.650 1531.940 1321.970 1532.000 ;
        RECT 1321.190 1531.800 1321.970 1531.940 ;
        RECT 1321.190 1531.740 1321.510 1531.800 ;
        RECT 1321.650 1531.740 1321.970 1531.800 ;
        RECT 1321.190 1483.660 1321.510 1483.720 ;
        RECT 1322.110 1483.660 1322.430 1483.720 ;
        RECT 1321.190 1483.520 1322.430 1483.660 ;
        RECT 1321.190 1483.460 1321.510 1483.520 ;
        RECT 1322.110 1483.460 1322.430 1483.520 ;
        RECT 1321.190 1186.840 1321.510 1186.900 ;
        RECT 1320.995 1186.700 1321.510 1186.840 ;
        RECT 1321.190 1186.640 1321.510 1186.700 ;
        RECT 1321.190 1097.420 1321.510 1097.480 ;
        RECT 1320.995 1097.280 1321.510 1097.420 ;
        RECT 1321.190 1097.220 1321.510 1097.280 ;
        RECT 1321.190 1089.940 1321.510 1090.000 ;
        RECT 1320.995 1089.800 1321.510 1089.940 ;
        RECT 1321.190 1089.740 1321.510 1089.800 ;
        RECT 1321.205 1042.000 1321.495 1042.045 ;
        RECT 1322.110 1042.000 1322.430 1042.060 ;
        RECT 1321.205 1041.860 1322.430 1042.000 ;
        RECT 1321.205 1041.815 1321.495 1041.860 ;
        RECT 1322.110 1041.800 1322.430 1041.860 ;
        RECT 1321.190 993.720 1321.510 993.780 ;
        RECT 1322.110 993.720 1322.430 993.780 ;
        RECT 1321.190 993.580 1322.430 993.720 ;
        RECT 1321.190 993.520 1321.510 993.580 ;
        RECT 1322.110 993.520 1322.430 993.580 ;
        RECT 1321.190 945.100 1321.510 945.160 ;
        RECT 1320.995 944.960 1321.510 945.100 ;
        RECT 1321.190 944.900 1321.510 944.960 ;
        RECT 1321.190 897.160 1321.510 897.220 ;
        RECT 1320.995 897.020 1321.510 897.160 ;
        RECT 1321.190 896.960 1321.510 897.020 ;
        RECT 1321.190 848.540 1321.510 848.600 ;
        RECT 1320.995 848.400 1321.510 848.540 ;
        RECT 1321.190 848.340 1321.510 848.400 ;
        RECT 1321.190 800.600 1321.510 800.660 ;
        RECT 1320.995 800.460 1321.510 800.600 ;
        RECT 1321.190 800.400 1321.510 800.460 ;
        RECT 1321.190 703.700 1321.510 703.760 ;
        RECT 1320.995 703.560 1321.510 703.700 ;
        RECT 1321.190 703.500 1321.510 703.560 ;
        RECT 1321.190 655.760 1321.510 655.820 ;
        RECT 1320.995 655.620 1321.510 655.760 ;
        RECT 1321.190 655.560 1321.510 655.620 ;
        RECT 1321.190 510.580 1321.510 510.640 ;
        RECT 1320.995 510.440 1321.510 510.580 ;
        RECT 1321.190 510.380 1321.510 510.440 ;
        RECT 1321.190 462.640 1321.510 462.700 ;
        RECT 1320.995 462.500 1321.510 462.640 ;
        RECT 1321.190 462.440 1321.510 462.500 ;
        RECT 1321.190 414.020 1321.510 414.080 ;
        RECT 1320.995 413.880 1321.510 414.020 ;
        RECT 1321.190 413.820 1321.510 413.880 ;
        RECT 1321.205 379.000 1321.495 379.045 ;
        RECT 1321.650 379.000 1321.970 379.060 ;
        RECT 1321.205 378.860 1321.970 379.000 ;
        RECT 1321.205 378.815 1321.495 378.860 ;
        RECT 1321.650 378.800 1321.970 378.860 ;
        RECT 1321.190 331.400 1321.510 331.460 ;
        RECT 1321.650 331.400 1321.970 331.460 ;
        RECT 1321.190 331.260 1321.970 331.400 ;
        RECT 1321.190 331.200 1321.510 331.260 ;
        RECT 1321.650 331.200 1321.970 331.260 ;
        RECT 1321.190 227.700 1321.510 227.760 ;
        RECT 1320.995 227.560 1321.510 227.700 ;
        RECT 1321.190 227.500 1321.510 227.560 ;
        RECT 1321.190 179.760 1321.510 179.820 ;
        RECT 1320.995 179.620 1321.510 179.760 ;
        RECT 1321.190 179.560 1321.510 179.620 ;
        RECT 1321.190 131.140 1321.510 131.200 ;
        RECT 1320.995 131.000 1321.510 131.140 ;
        RECT 1321.190 130.940 1321.510 131.000 ;
        RECT 1321.190 83.200 1321.510 83.260 ;
        RECT 1320.995 83.060 1321.510 83.200 ;
        RECT 1321.190 83.000 1321.510 83.060 ;
        RECT 1321.190 34.240 1321.510 34.300 ;
        RECT 1320.995 34.100 1321.510 34.240 ;
        RECT 1321.190 34.040 1321.510 34.100 ;
        RECT 1321.205 28.460 1321.495 28.505 ;
        RECT 1650.090 28.460 1650.410 28.520 ;
        RECT 1321.205 28.320 1650.410 28.460 ;
        RECT 1321.205 28.275 1321.495 28.320 ;
        RECT 1650.090 28.260 1650.410 28.320 ;
      LAYER via ;
        RECT 1319.380 1634.760 1319.640 1635.020 ;
        RECT 1321.680 1634.760 1321.940 1635.020 ;
        RECT 1321.220 1531.740 1321.480 1532.000 ;
        RECT 1321.680 1531.740 1321.940 1532.000 ;
        RECT 1321.220 1483.460 1321.480 1483.720 ;
        RECT 1322.140 1483.460 1322.400 1483.720 ;
        RECT 1321.220 1186.640 1321.480 1186.900 ;
        RECT 1321.220 1097.220 1321.480 1097.480 ;
        RECT 1321.220 1089.740 1321.480 1090.000 ;
        RECT 1322.140 1041.800 1322.400 1042.060 ;
        RECT 1321.220 993.520 1321.480 993.780 ;
        RECT 1322.140 993.520 1322.400 993.780 ;
        RECT 1321.220 944.900 1321.480 945.160 ;
        RECT 1321.220 896.960 1321.480 897.220 ;
        RECT 1321.220 848.340 1321.480 848.600 ;
        RECT 1321.220 800.400 1321.480 800.660 ;
        RECT 1321.220 703.500 1321.480 703.760 ;
        RECT 1321.220 655.560 1321.480 655.820 ;
        RECT 1321.220 510.380 1321.480 510.640 ;
        RECT 1321.220 462.440 1321.480 462.700 ;
        RECT 1321.220 413.820 1321.480 414.080 ;
        RECT 1321.680 378.800 1321.940 379.060 ;
        RECT 1321.220 331.200 1321.480 331.460 ;
        RECT 1321.680 331.200 1321.940 331.460 ;
        RECT 1321.220 227.500 1321.480 227.760 ;
        RECT 1321.220 179.560 1321.480 179.820 ;
        RECT 1321.220 130.940 1321.480 131.200 ;
        RECT 1321.220 83.000 1321.480 83.260 ;
        RECT 1321.220 34.040 1321.480 34.300 ;
        RECT 1650.120 28.260 1650.380 28.520 ;
      LAYER met2 ;
        RECT 1319.280 1700.340 1319.560 1704.000 ;
        RECT 1319.280 1700.000 1319.580 1700.340 ;
        RECT 1319.440 1635.050 1319.580 1700.000 ;
        RECT 1319.380 1634.730 1319.640 1635.050 ;
        RECT 1321.680 1634.730 1321.940 1635.050 ;
        RECT 1321.740 1532.030 1321.880 1634.730 ;
        RECT 1321.220 1531.885 1321.480 1532.030 ;
        RECT 1321.210 1531.515 1321.490 1531.885 ;
        RECT 1321.680 1531.710 1321.940 1532.030 ;
        RECT 1322.130 1531.515 1322.410 1531.885 ;
        RECT 1322.200 1483.750 1322.340 1531.515 ;
        RECT 1321.220 1483.430 1321.480 1483.750 ;
        RECT 1322.140 1483.430 1322.400 1483.750 ;
        RECT 1321.280 1186.930 1321.420 1483.430 ;
        RECT 1321.220 1186.610 1321.480 1186.930 ;
        RECT 1321.220 1097.190 1321.480 1097.510 ;
        RECT 1321.280 1090.030 1321.420 1097.190 ;
        RECT 1321.220 1089.710 1321.480 1090.030 ;
        RECT 1322.140 1041.770 1322.400 1042.090 ;
        RECT 1322.200 993.810 1322.340 1041.770 ;
        RECT 1321.220 993.490 1321.480 993.810 ;
        RECT 1322.140 993.490 1322.400 993.810 ;
        RECT 1321.280 945.190 1321.420 993.490 ;
        RECT 1321.220 944.870 1321.480 945.190 ;
        RECT 1321.220 896.930 1321.480 897.250 ;
        RECT 1321.280 848.630 1321.420 896.930 ;
        RECT 1321.220 848.310 1321.480 848.630 ;
        RECT 1321.220 800.370 1321.480 800.690 ;
        RECT 1321.280 703.790 1321.420 800.370 ;
        RECT 1321.220 703.470 1321.480 703.790 ;
        RECT 1321.220 655.530 1321.480 655.850 ;
        RECT 1321.280 510.670 1321.420 655.530 ;
        RECT 1321.220 510.350 1321.480 510.670 ;
        RECT 1321.220 462.410 1321.480 462.730 ;
        RECT 1321.280 462.130 1321.420 462.410 ;
        RECT 1321.280 461.990 1321.880 462.130 ;
        RECT 1321.740 414.530 1321.880 461.990 ;
        RECT 1321.280 414.390 1321.880 414.530 ;
        RECT 1321.280 414.110 1321.420 414.390 ;
        RECT 1321.220 413.790 1321.480 414.110 ;
        RECT 1321.680 378.770 1321.940 379.090 ;
        RECT 1321.740 331.490 1321.880 378.770 ;
        RECT 1321.220 331.170 1321.480 331.490 ;
        RECT 1321.680 331.170 1321.940 331.490 ;
        RECT 1321.280 227.790 1321.420 331.170 ;
        RECT 1321.220 227.470 1321.480 227.790 ;
        RECT 1321.220 179.530 1321.480 179.850 ;
        RECT 1321.280 131.230 1321.420 179.530 ;
        RECT 1321.220 130.910 1321.480 131.230 ;
        RECT 1321.220 82.970 1321.480 83.290 ;
        RECT 1321.280 34.330 1321.420 82.970 ;
        RECT 1321.220 34.010 1321.480 34.330 ;
        RECT 1650.120 28.230 1650.380 28.550 ;
        RECT 1650.180 2.400 1650.320 28.230 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
      LAYER via2 ;
        RECT 1321.210 1531.560 1321.490 1531.840 ;
        RECT 1322.130 1531.560 1322.410 1531.840 ;
      LAYER met3 ;
        RECT 1321.185 1531.850 1321.515 1531.865 ;
        RECT 1322.105 1531.850 1322.435 1531.865 ;
        RECT 1321.185 1531.550 1322.435 1531.850 ;
        RECT 1321.185 1531.535 1321.515 1531.550 ;
        RECT 1322.105 1531.535 1322.435 1531.550 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1320.270 1631.900 1320.590 1631.960 ;
        RECT 1321.190 1631.900 1321.510 1631.960 ;
        RECT 1320.270 1631.760 1321.510 1631.900 ;
        RECT 1320.270 1631.700 1320.590 1631.760 ;
        RECT 1321.190 1631.700 1321.510 1631.760 ;
        RECT 1320.270 28.800 1320.590 28.860 ;
        RECT 1668.030 28.800 1668.350 28.860 ;
        RECT 1320.270 28.660 1668.350 28.800 ;
        RECT 1320.270 28.600 1320.590 28.660 ;
        RECT 1668.030 28.600 1668.350 28.660 ;
      LAYER via ;
        RECT 1320.300 1631.700 1320.560 1631.960 ;
        RECT 1321.220 1631.700 1321.480 1631.960 ;
        RECT 1320.300 28.600 1320.560 28.860 ;
        RECT 1668.060 28.600 1668.320 28.860 ;
      LAYER met2 ;
        RECT 1321.120 1700.340 1321.400 1704.000 ;
        RECT 1321.120 1700.000 1321.420 1700.340 ;
        RECT 1321.280 1631.990 1321.420 1700.000 ;
        RECT 1320.300 1631.670 1320.560 1631.990 ;
        RECT 1321.220 1631.670 1321.480 1631.990 ;
        RECT 1320.360 28.890 1320.500 1631.670 ;
        RECT 1320.300 28.570 1320.560 28.890 ;
        RECT 1668.060 28.570 1668.320 28.890 ;
        RECT 1668.120 2.400 1668.260 28.570 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1320.730 1684.260 1321.050 1684.320 ;
        RECT 1323.030 1684.260 1323.350 1684.320 ;
        RECT 1320.730 1684.120 1323.350 1684.260 ;
        RECT 1320.730 1684.060 1321.050 1684.120 ;
        RECT 1323.030 1684.060 1323.350 1684.120 ;
        RECT 1320.730 29.140 1321.050 29.200 ;
        RECT 1685.510 29.140 1685.830 29.200 ;
        RECT 1320.730 29.000 1685.830 29.140 ;
        RECT 1320.730 28.940 1321.050 29.000 ;
        RECT 1685.510 28.940 1685.830 29.000 ;
      LAYER via ;
        RECT 1320.760 1684.060 1321.020 1684.320 ;
        RECT 1323.060 1684.060 1323.320 1684.320 ;
        RECT 1320.760 28.940 1321.020 29.200 ;
        RECT 1685.540 28.940 1685.800 29.200 ;
      LAYER met2 ;
        RECT 1322.960 1700.340 1323.240 1704.000 ;
        RECT 1322.960 1700.000 1323.260 1700.340 ;
        RECT 1323.120 1684.350 1323.260 1700.000 ;
        RECT 1320.760 1684.030 1321.020 1684.350 ;
        RECT 1323.060 1684.030 1323.320 1684.350 ;
        RECT 1320.820 29.230 1320.960 1684.030 ;
        RECT 1320.760 28.910 1321.020 29.230 ;
        RECT 1685.540 28.910 1685.800 29.230 ;
        RECT 1685.600 2.400 1685.740 28.910 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1224.130 1678.480 1224.450 1678.540 ;
        RECT 1225.510 1678.480 1225.830 1678.540 ;
        RECT 1224.130 1678.340 1225.830 1678.480 ;
        RECT 1224.130 1678.280 1224.450 1678.340 ;
        RECT 1225.510 1678.280 1225.830 1678.340 ;
        RECT 724.110 1660.120 724.430 1660.180 ;
        RECT 1225.510 1660.120 1225.830 1660.180 ;
        RECT 724.110 1659.980 1225.830 1660.120 ;
        RECT 724.110 1659.920 724.430 1659.980 ;
        RECT 1225.510 1659.920 1225.830 1659.980 ;
      LAYER via ;
        RECT 1224.160 1678.280 1224.420 1678.540 ;
        RECT 1225.540 1678.280 1225.800 1678.540 ;
        RECT 724.140 1659.920 724.400 1660.180 ;
        RECT 1225.540 1659.920 1225.800 1660.180 ;
      LAYER met2 ;
        RECT 1224.060 1700.340 1224.340 1704.000 ;
        RECT 1224.060 1700.000 1224.360 1700.340 ;
        RECT 1224.220 1678.570 1224.360 1700.000 ;
        RECT 1224.160 1678.250 1224.420 1678.570 ;
        RECT 1225.540 1678.250 1225.800 1678.570 ;
        RECT 1225.600 1660.210 1225.740 1678.250 ;
        RECT 724.140 1659.890 724.400 1660.210 ;
        RECT 1225.540 1659.890 1225.800 1660.210 ;
        RECT 724.200 16.730 724.340 1659.890 ;
        RECT 722.360 16.590 724.340 16.730 ;
        RECT 722.360 2.400 722.500 16.590 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1324.870 29.480 1325.190 29.540 ;
        RECT 1703.450 29.480 1703.770 29.540 ;
        RECT 1324.870 29.340 1703.770 29.480 ;
        RECT 1324.870 29.280 1325.190 29.340 ;
        RECT 1703.450 29.280 1703.770 29.340 ;
      LAYER via ;
        RECT 1324.900 29.280 1325.160 29.540 ;
        RECT 1703.480 29.280 1703.740 29.540 ;
      LAYER met2 ;
        RECT 1324.800 1700.340 1325.080 1704.000 ;
        RECT 1324.800 1700.000 1325.100 1700.340 ;
        RECT 1324.960 29.570 1325.100 1700.000 ;
        RECT 1324.900 29.250 1325.160 29.570 ;
        RECT 1703.480 29.250 1703.740 29.570 ;
        RECT 1703.540 2.400 1703.680 29.250 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1331.385 1635.485 1331.555 1683.595 ;
      LAYER mcon ;
        RECT 1331.385 1683.425 1331.555 1683.595 ;
      LAYER met1 ;
        RECT 1326.710 1684.260 1327.030 1684.320 ;
        RECT 1331.310 1684.260 1331.630 1684.320 ;
        RECT 1326.710 1684.120 1331.630 1684.260 ;
        RECT 1326.710 1684.060 1327.030 1684.120 ;
        RECT 1331.310 1684.060 1331.630 1684.120 ;
        RECT 1331.310 1683.580 1331.630 1683.640 ;
        RECT 1331.115 1683.440 1331.630 1683.580 ;
        RECT 1331.310 1683.380 1331.630 1683.440 ;
        RECT 1331.310 1635.640 1331.630 1635.700 ;
        RECT 1331.115 1635.500 1331.630 1635.640 ;
        RECT 1331.310 1635.440 1331.630 1635.500 ;
        RECT 1330.850 1497.600 1331.170 1497.660 ;
        RECT 1331.310 1497.600 1331.630 1497.660 ;
        RECT 1330.850 1497.460 1331.630 1497.600 ;
        RECT 1330.850 1497.400 1331.170 1497.460 ;
        RECT 1331.310 1497.400 1331.630 1497.460 ;
        RECT 1330.850 29.820 1331.170 29.880 ;
        RECT 1721.390 29.820 1721.710 29.880 ;
        RECT 1330.850 29.680 1721.710 29.820 ;
        RECT 1330.850 29.620 1331.170 29.680 ;
        RECT 1721.390 29.620 1721.710 29.680 ;
      LAYER via ;
        RECT 1326.740 1684.060 1327.000 1684.320 ;
        RECT 1331.340 1684.060 1331.600 1684.320 ;
        RECT 1331.340 1683.380 1331.600 1683.640 ;
        RECT 1331.340 1635.440 1331.600 1635.700 ;
        RECT 1330.880 1497.400 1331.140 1497.660 ;
        RECT 1331.340 1497.400 1331.600 1497.660 ;
        RECT 1330.880 29.620 1331.140 29.880 ;
        RECT 1721.420 29.620 1721.680 29.880 ;
      LAYER met2 ;
        RECT 1326.640 1700.340 1326.920 1704.000 ;
        RECT 1326.640 1700.000 1326.940 1700.340 ;
        RECT 1326.800 1684.350 1326.940 1700.000 ;
        RECT 1326.740 1684.030 1327.000 1684.350 ;
        RECT 1331.340 1684.030 1331.600 1684.350 ;
        RECT 1331.400 1683.670 1331.540 1684.030 ;
        RECT 1331.340 1683.350 1331.600 1683.670 ;
        RECT 1331.340 1635.410 1331.600 1635.730 ;
        RECT 1331.400 1497.690 1331.540 1635.410 ;
        RECT 1330.880 1497.370 1331.140 1497.690 ;
        RECT 1331.340 1497.370 1331.600 1497.690 ;
        RECT 1330.940 29.910 1331.080 1497.370 ;
        RECT 1330.880 29.590 1331.140 29.910 ;
        RECT 1721.420 29.590 1721.680 29.910 ;
        RECT 1721.480 2.400 1721.620 29.590 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1328.550 1677.460 1328.870 1677.520 ;
        RECT 1330.390 1677.460 1330.710 1677.520 ;
        RECT 1328.550 1677.320 1330.710 1677.460 ;
        RECT 1328.550 1677.260 1328.870 1677.320 ;
        RECT 1330.390 1677.260 1330.710 1677.320 ;
        RECT 1330.390 30.160 1330.710 30.220 ;
        RECT 1739.330 30.160 1739.650 30.220 ;
        RECT 1330.390 30.020 1739.650 30.160 ;
        RECT 1330.390 29.960 1330.710 30.020 ;
        RECT 1739.330 29.960 1739.650 30.020 ;
      LAYER via ;
        RECT 1328.580 1677.260 1328.840 1677.520 ;
        RECT 1330.420 1677.260 1330.680 1677.520 ;
        RECT 1330.420 29.960 1330.680 30.220 ;
        RECT 1739.360 29.960 1739.620 30.220 ;
      LAYER met2 ;
        RECT 1328.480 1700.340 1328.760 1704.000 ;
        RECT 1328.480 1700.000 1328.780 1700.340 ;
        RECT 1328.640 1677.550 1328.780 1700.000 ;
        RECT 1328.580 1677.230 1328.840 1677.550 ;
        RECT 1330.420 1677.230 1330.680 1677.550 ;
        RECT 1330.480 30.250 1330.620 1677.230 ;
        RECT 1330.420 29.930 1330.680 30.250 ;
        RECT 1739.360 29.930 1739.620 30.250 ;
        RECT 1739.420 2.400 1739.560 29.930 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1327.245 1636.845 1327.415 1678.495 ;
      LAYER mcon ;
        RECT 1327.245 1678.325 1327.415 1678.495 ;
      LAYER met1 ;
        RECT 1327.185 1678.480 1327.475 1678.525 ;
        RECT 1330.390 1678.480 1330.710 1678.540 ;
        RECT 1327.185 1678.340 1330.710 1678.480 ;
        RECT 1327.185 1678.295 1327.475 1678.340 ;
        RECT 1330.390 1678.280 1330.710 1678.340 ;
        RECT 1327.170 1637.000 1327.490 1637.060 ;
        RECT 1326.975 1636.860 1327.490 1637.000 ;
        RECT 1327.170 1636.800 1327.490 1636.860 ;
        RECT 1327.170 30.500 1327.490 30.560 ;
        RECT 1756.810 30.500 1757.130 30.560 ;
        RECT 1327.170 30.360 1757.130 30.500 ;
        RECT 1327.170 30.300 1327.490 30.360 ;
        RECT 1756.810 30.300 1757.130 30.360 ;
      LAYER via ;
        RECT 1330.420 1678.280 1330.680 1678.540 ;
        RECT 1327.200 1636.800 1327.460 1637.060 ;
        RECT 1327.200 30.300 1327.460 30.560 ;
        RECT 1756.840 30.300 1757.100 30.560 ;
      LAYER met2 ;
        RECT 1330.320 1700.340 1330.600 1704.000 ;
        RECT 1330.320 1700.000 1330.620 1700.340 ;
        RECT 1330.480 1678.570 1330.620 1700.000 ;
        RECT 1330.420 1678.250 1330.680 1678.570 ;
        RECT 1327.200 1636.770 1327.460 1637.090 ;
        RECT 1327.260 30.590 1327.400 1636.770 ;
        RECT 1327.200 30.270 1327.460 30.590 ;
        RECT 1756.840 30.270 1757.100 30.590 ;
        RECT 1756.900 2.400 1757.040 30.270 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1333.150 1631.900 1333.470 1631.960 ;
        RECT 1334.070 1631.900 1334.390 1631.960 ;
        RECT 1333.150 1631.760 1334.390 1631.900 ;
        RECT 1333.150 1631.700 1333.470 1631.760 ;
        RECT 1334.070 1631.700 1334.390 1631.760 ;
        RECT 1334.070 34.240 1334.390 34.300 ;
        RECT 1774.750 34.240 1775.070 34.300 ;
        RECT 1334.070 34.100 1775.070 34.240 ;
        RECT 1334.070 34.040 1334.390 34.100 ;
        RECT 1774.750 34.040 1775.070 34.100 ;
      LAYER via ;
        RECT 1333.180 1631.700 1333.440 1631.960 ;
        RECT 1334.100 1631.700 1334.360 1631.960 ;
        RECT 1334.100 34.040 1334.360 34.300 ;
        RECT 1774.780 34.040 1775.040 34.300 ;
      LAYER met2 ;
        RECT 1332.160 1700.340 1332.440 1704.000 ;
        RECT 1332.160 1700.000 1332.460 1700.340 ;
        RECT 1332.320 1677.970 1332.460 1700.000 ;
        RECT 1332.320 1677.830 1333.380 1677.970 ;
        RECT 1333.240 1631.990 1333.380 1677.830 ;
        RECT 1333.180 1631.670 1333.440 1631.990 ;
        RECT 1334.100 1631.670 1334.360 1631.990 ;
        RECT 1334.160 34.330 1334.300 1631.670 ;
        RECT 1334.100 34.010 1334.360 34.330 ;
        RECT 1774.780 34.010 1775.040 34.330 ;
        RECT 1774.840 2.400 1774.980 34.010 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1333.610 33.900 1333.930 33.960 ;
        RECT 1792.690 33.900 1793.010 33.960 ;
        RECT 1333.610 33.760 1793.010 33.900 ;
        RECT 1333.610 33.700 1333.930 33.760 ;
        RECT 1792.690 33.700 1793.010 33.760 ;
      LAYER via ;
        RECT 1333.640 33.700 1333.900 33.960 ;
        RECT 1792.720 33.700 1792.980 33.960 ;
      LAYER met2 ;
        RECT 1334.000 1700.340 1334.280 1704.000 ;
        RECT 1334.000 1700.000 1334.300 1700.340 ;
        RECT 1334.160 1659.610 1334.300 1700.000 ;
        RECT 1333.700 1659.470 1334.300 1659.610 ;
        RECT 1333.700 33.990 1333.840 1659.470 ;
        RECT 1333.640 33.670 1333.900 33.990 ;
        RECT 1792.720 33.670 1792.980 33.990 ;
        RECT 1792.780 2.400 1792.920 33.670 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1331.770 1684.940 1332.090 1685.000 ;
        RECT 1335.910 1684.940 1336.230 1685.000 ;
        RECT 1331.770 1684.800 1336.230 1684.940 ;
        RECT 1331.770 1684.740 1332.090 1684.800 ;
        RECT 1335.910 1684.740 1336.230 1684.800 ;
        RECT 1332.690 33.560 1333.010 33.620 ;
        RECT 1810.630 33.560 1810.950 33.620 ;
        RECT 1332.690 33.420 1810.950 33.560 ;
        RECT 1332.690 33.360 1333.010 33.420 ;
        RECT 1810.630 33.360 1810.950 33.420 ;
      LAYER via ;
        RECT 1331.800 1684.740 1332.060 1685.000 ;
        RECT 1335.940 1684.740 1336.200 1685.000 ;
        RECT 1332.720 33.360 1332.980 33.620 ;
        RECT 1810.660 33.360 1810.920 33.620 ;
      LAYER met2 ;
        RECT 1335.840 1700.340 1336.120 1704.000 ;
        RECT 1335.840 1700.000 1336.140 1700.340 ;
        RECT 1336.000 1685.030 1336.140 1700.000 ;
        RECT 1331.800 1684.710 1332.060 1685.030 ;
        RECT 1335.940 1684.710 1336.200 1685.030 ;
        RECT 1331.860 1677.290 1332.000 1684.710 ;
        RECT 1331.860 1677.150 1332.920 1677.290 ;
        RECT 1332.780 33.650 1332.920 1677.150 ;
        RECT 1332.720 33.330 1332.980 33.650 ;
        RECT 1810.660 33.330 1810.920 33.650 ;
        RECT 1810.720 2.400 1810.860 33.330 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1333.610 1686.300 1333.930 1686.360 ;
        RECT 1337.750 1686.300 1338.070 1686.360 ;
        RECT 1333.610 1686.160 1338.070 1686.300 ;
        RECT 1333.610 1686.100 1333.930 1686.160 ;
        RECT 1337.750 1686.100 1338.070 1686.160 ;
        RECT 1332.230 1660.120 1332.550 1660.180 ;
        RECT 1333.610 1660.120 1333.930 1660.180 ;
        RECT 1332.230 1659.980 1333.930 1660.120 ;
        RECT 1332.230 1659.920 1332.550 1659.980 ;
        RECT 1333.610 1659.920 1333.930 1659.980 ;
        RECT 1332.230 33.220 1332.550 33.280 ;
        RECT 1829.030 33.220 1829.350 33.280 ;
        RECT 1332.230 33.080 1829.350 33.220 ;
        RECT 1332.230 33.020 1332.550 33.080 ;
        RECT 1829.030 33.020 1829.350 33.080 ;
      LAYER via ;
        RECT 1333.640 1686.100 1333.900 1686.360 ;
        RECT 1337.780 1686.100 1338.040 1686.360 ;
        RECT 1332.260 1659.920 1332.520 1660.180 ;
        RECT 1333.640 1659.920 1333.900 1660.180 ;
        RECT 1332.260 33.020 1332.520 33.280 ;
        RECT 1829.060 33.020 1829.320 33.280 ;
      LAYER met2 ;
        RECT 1337.680 1700.340 1337.960 1704.000 ;
        RECT 1337.680 1700.000 1337.980 1700.340 ;
        RECT 1337.840 1686.390 1337.980 1700.000 ;
        RECT 1333.640 1686.070 1333.900 1686.390 ;
        RECT 1337.780 1686.070 1338.040 1686.390 ;
        RECT 1333.700 1660.210 1333.840 1686.070 ;
        RECT 1332.260 1659.890 1332.520 1660.210 ;
        RECT 1333.640 1659.890 1333.900 1660.210 ;
        RECT 1332.320 33.310 1332.460 1659.890 ;
        RECT 1332.260 32.990 1332.520 33.310 ;
        RECT 1829.060 32.990 1829.320 33.310 ;
        RECT 1829.120 16.730 1829.260 32.990 ;
        RECT 1828.660 16.590 1829.260 16.730 ;
        RECT 1828.660 2.400 1828.800 16.590 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1341.430 32.880 1341.750 32.940 ;
        RECT 1846.050 32.880 1846.370 32.940 ;
        RECT 1341.430 32.740 1846.370 32.880 ;
        RECT 1341.430 32.680 1341.750 32.740 ;
        RECT 1846.050 32.680 1846.370 32.740 ;
      LAYER via ;
        RECT 1341.460 32.680 1341.720 32.940 ;
        RECT 1846.080 32.680 1846.340 32.940 ;
      LAYER met2 ;
        RECT 1339.520 1700.340 1339.800 1704.000 ;
        RECT 1339.520 1700.000 1339.820 1700.340 ;
        RECT 1339.680 1677.970 1339.820 1700.000 ;
        RECT 1339.680 1677.830 1340.740 1677.970 ;
        RECT 1340.600 169.050 1340.740 1677.830 ;
        RECT 1340.600 168.910 1341.660 169.050 ;
        RECT 1341.520 32.970 1341.660 168.910 ;
        RECT 1341.460 32.650 1341.720 32.970 ;
        RECT 1846.080 32.650 1846.340 32.970 ;
        RECT 1846.140 2.400 1846.280 32.650 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1338.670 1683.920 1338.990 1683.980 ;
        RECT 1341.430 1683.920 1341.750 1683.980 ;
        RECT 1338.670 1683.780 1341.750 1683.920 ;
        RECT 1338.670 1683.720 1338.990 1683.780 ;
        RECT 1341.430 1683.720 1341.750 1683.780 ;
        RECT 1338.670 1631.900 1338.990 1631.960 ;
        RECT 1339.590 1631.900 1339.910 1631.960 ;
        RECT 1338.670 1631.760 1339.910 1631.900 ;
        RECT 1338.670 1631.700 1338.990 1631.760 ;
        RECT 1339.590 1631.700 1339.910 1631.760 ;
        RECT 1339.590 32.540 1339.910 32.600 ;
        RECT 1863.990 32.540 1864.310 32.600 ;
        RECT 1339.590 32.400 1864.310 32.540 ;
        RECT 1339.590 32.340 1339.910 32.400 ;
        RECT 1863.990 32.340 1864.310 32.400 ;
      LAYER via ;
        RECT 1338.700 1683.720 1338.960 1683.980 ;
        RECT 1341.460 1683.720 1341.720 1683.980 ;
        RECT 1338.700 1631.700 1338.960 1631.960 ;
        RECT 1339.620 1631.700 1339.880 1631.960 ;
        RECT 1339.620 32.340 1339.880 32.600 ;
        RECT 1864.020 32.340 1864.280 32.600 ;
      LAYER met2 ;
        RECT 1341.360 1700.340 1341.640 1704.000 ;
        RECT 1341.360 1700.000 1341.660 1700.340 ;
        RECT 1341.520 1684.010 1341.660 1700.000 ;
        RECT 1338.700 1683.690 1338.960 1684.010 ;
        RECT 1341.460 1683.690 1341.720 1684.010 ;
        RECT 1338.760 1631.990 1338.900 1683.690 ;
        RECT 1338.700 1631.670 1338.960 1631.990 ;
        RECT 1339.620 1631.670 1339.880 1631.990 ;
        RECT 1339.680 32.630 1339.820 1631.670 ;
        RECT 1339.620 32.310 1339.880 32.630 ;
        RECT 1864.020 32.310 1864.280 32.630 ;
        RECT 1864.080 2.400 1864.220 32.310 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1128.450 1685.960 1128.770 1686.020 ;
        RECT 1225.510 1685.960 1225.830 1686.020 ;
        RECT 1128.450 1685.820 1225.830 1685.960 ;
        RECT 1128.450 1685.760 1128.770 1685.820 ;
        RECT 1225.510 1685.760 1225.830 1685.820 ;
        RECT 744.810 65.520 745.130 65.580 ;
        RECT 1128.450 65.520 1128.770 65.580 ;
        RECT 744.810 65.380 1128.770 65.520 ;
        RECT 744.810 65.320 745.130 65.380 ;
        RECT 1128.450 65.320 1128.770 65.380 ;
      LAYER via ;
        RECT 1128.480 1685.760 1128.740 1686.020 ;
        RECT 1225.540 1685.760 1225.800 1686.020 ;
        RECT 744.840 65.320 745.100 65.580 ;
        RECT 1128.480 65.320 1128.740 65.580 ;
      LAYER met2 ;
        RECT 1225.440 1700.340 1225.720 1704.000 ;
        RECT 1225.440 1700.000 1225.740 1700.340 ;
        RECT 1225.600 1686.050 1225.740 1700.000 ;
        RECT 1128.480 1685.730 1128.740 1686.050 ;
        RECT 1225.540 1685.730 1225.800 1686.050 ;
        RECT 1128.540 65.610 1128.680 1685.730 ;
        RECT 744.840 65.290 745.100 65.610 ;
        RECT 1128.480 65.290 1128.740 65.610 ;
        RECT 744.900 16.730 745.040 65.290 ;
        RECT 740.300 16.590 745.040 16.730 ;
        RECT 740.300 2.400 740.440 16.590 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1340.050 1685.960 1340.370 1686.020 ;
        RECT 1343.270 1685.960 1343.590 1686.020 ;
        RECT 1340.050 1685.820 1343.590 1685.960 ;
        RECT 1340.050 1685.760 1340.370 1685.820 ;
        RECT 1343.270 1685.760 1343.590 1685.820 ;
        RECT 1340.050 1678.280 1340.370 1678.540 ;
        RECT 1340.140 1677.520 1340.280 1678.280 ;
        RECT 1340.050 1677.260 1340.370 1677.520 ;
        RECT 1340.050 32.200 1340.370 32.260 ;
        RECT 1881.930 32.200 1882.250 32.260 ;
        RECT 1340.050 32.060 1882.250 32.200 ;
        RECT 1340.050 32.000 1340.370 32.060 ;
        RECT 1881.930 32.000 1882.250 32.060 ;
      LAYER via ;
        RECT 1340.080 1685.760 1340.340 1686.020 ;
        RECT 1343.300 1685.760 1343.560 1686.020 ;
        RECT 1340.080 1678.280 1340.340 1678.540 ;
        RECT 1340.080 1677.260 1340.340 1677.520 ;
        RECT 1340.080 32.000 1340.340 32.260 ;
        RECT 1881.960 32.000 1882.220 32.260 ;
      LAYER met2 ;
        RECT 1343.200 1700.340 1343.480 1704.000 ;
        RECT 1343.200 1700.000 1343.500 1700.340 ;
        RECT 1343.360 1686.050 1343.500 1700.000 ;
        RECT 1340.080 1685.730 1340.340 1686.050 ;
        RECT 1343.300 1685.730 1343.560 1686.050 ;
        RECT 1340.140 1678.570 1340.280 1685.730 ;
        RECT 1340.080 1678.250 1340.340 1678.570 ;
        RECT 1340.080 1677.230 1340.340 1677.550 ;
        RECT 1340.140 32.290 1340.280 1677.230 ;
        RECT 1340.080 31.970 1340.340 32.290 ;
        RECT 1881.960 31.970 1882.220 32.290 ;
        RECT 1882.020 2.400 1882.160 31.970 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1344.650 1683.920 1344.970 1683.980 ;
        RECT 1341.980 1683.780 1344.970 1683.920 ;
        RECT 1339.130 1683.580 1339.450 1683.640 ;
        RECT 1341.980 1683.580 1342.120 1683.780 ;
        RECT 1344.650 1683.720 1344.970 1683.780 ;
        RECT 1339.130 1683.440 1342.120 1683.580 ;
        RECT 1339.130 1683.380 1339.450 1683.440 ;
        RECT 1339.130 31.860 1339.450 31.920 ;
        RECT 1899.870 31.860 1900.190 31.920 ;
        RECT 1339.130 31.720 1900.190 31.860 ;
        RECT 1339.130 31.660 1339.450 31.720 ;
        RECT 1899.870 31.660 1900.190 31.720 ;
      LAYER via ;
        RECT 1339.160 1683.380 1339.420 1683.640 ;
        RECT 1344.680 1683.720 1344.940 1683.980 ;
        RECT 1339.160 31.660 1339.420 31.920 ;
        RECT 1899.900 31.660 1900.160 31.920 ;
      LAYER met2 ;
        RECT 1345.040 1700.340 1345.320 1704.000 ;
        RECT 1345.040 1700.000 1345.340 1700.340 ;
        RECT 1345.200 1687.490 1345.340 1700.000 ;
        RECT 1344.740 1687.350 1345.340 1687.490 ;
        RECT 1344.740 1684.010 1344.880 1687.350 ;
        RECT 1344.680 1683.690 1344.940 1684.010 ;
        RECT 1339.160 1683.350 1339.420 1683.670 ;
        RECT 1339.220 31.950 1339.360 1683.350 ;
        RECT 1339.160 31.630 1339.420 31.950 ;
        RECT 1899.900 31.630 1900.160 31.950 ;
        RECT 1899.960 2.400 1900.100 31.630 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.950 1684.940 1347.270 1685.000 ;
        RECT 1346.950 1684.800 1351.320 1684.940 ;
        RECT 1346.950 1684.740 1347.270 1684.800 ;
        RECT 1351.180 1683.920 1351.320 1684.800 ;
        RECT 1350.720 1683.780 1351.320 1683.920 ;
        RECT 1350.720 1683.640 1350.860 1683.780 ;
        RECT 1350.630 1683.380 1350.950 1683.640 ;
        RECT 1350.630 31.520 1350.950 31.580 ;
        RECT 1917.810 31.520 1918.130 31.580 ;
        RECT 1350.630 31.380 1918.130 31.520 ;
        RECT 1350.630 31.320 1350.950 31.380 ;
        RECT 1917.810 31.320 1918.130 31.380 ;
      LAYER via ;
        RECT 1346.980 1684.740 1347.240 1685.000 ;
        RECT 1350.660 1683.380 1350.920 1683.640 ;
        RECT 1350.660 31.320 1350.920 31.580 ;
        RECT 1917.840 31.320 1918.100 31.580 ;
      LAYER met2 ;
        RECT 1346.880 1700.340 1347.160 1704.000 ;
        RECT 1346.880 1700.000 1347.180 1700.340 ;
        RECT 1347.040 1685.030 1347.180 1700.000 ;
        RECT 1346.980 1684.710 1347.240 1685.030 ;
        RECT 1350.660 1683.350 1350.920 1683.670 ;
        RECT 1350.720 31.610 1350.860 1683.350 ;
        RECT 1350.660 31.290 1350.920 31.610 ;
        RECT 1917.840 31.290 1918.100 31.610 ;
        RECT 1917.900 2.400 1918.040 31.290 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.950 1683.920 1347.270 1683.980 ;
        RECT 1348.790 1683.920 1349.110 1683.980 ;
        RECT 1346.950 1683.780 1349.110 1683.920 ;
        RECT 1346.950 1683.720 1347.270 1683.780 ;
        RECT 1348.790 1683.720 1349.110 1683.780 ;
        RECT 1346.950 31.180 1347.270 31.240 ;
        RECT 1935.290 31.180 1935.610 31.240 ;
        RECT 1346.950 31.040 1935.610 31.180 ;
        RECT 1346.950 30.980 1347.270 31.040 ;
        RECT 1935.290 30.980 1935.610 31.040 ;
      LAYER via ;
        RECT 1346.980 1683.720 1347.240 1683.980 ;
        RECT 1348.820 1683.720 1349.080 1683.980 ;
        RECT 1346.980 30.980 1347.240 31.240 ;
        RECT 1935.320 30.980 1935.580 31.240 ;
      LAYER met2 ;
        RECT 1348.720 1700.340 1349.000 1704.000 ;
        RECT 1348.720 1700.000 1349.020 1700.340 ;
        RECT 1348.880 1684.010 1349.020 1700.000 ;
        RECT 1346.980 1683.690 1347.240 1684.010 ;
        RECT 1348.820 1683.690 1349.080 1684.010 ;
        RECT 1347.040 31.270 1347.180 1683.690 ;
        RECT 1346.980 30.950 1347.240 31.270 ;
        RECT 1935.320 30.950 1935.580 31.270 ;
        RECT 1935.380 2.400 1935.520 30.950 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1347.870 1684.260 1348.190 1684.320 ;
        RECT 1350.630 1684.260 1350.950 1684.320 ;
        RECT 1347.870 1684.120 1350.950 1684.260 ;
        RECT 1347.870 1684.060 1348.190 1684.120 ;
        RECT 1350.630 1684.060 1350.950 1684.120 ;
        RECT 1347.870 1634.760 1348.190 1635.020 ;
        RECT 1347.410 1633.940 1347.730 1634.000 ;
        RECT 1347.960 1633.940 1348.100 1634.760 ;
        RECT 1347.410 1633.800 1348.100 1633.940 ;
        RECT 1347.410 1633.740 1347.730 1633.800 ;
        RECT 1347.410 30.840 1347.730 30.900 ;
        RECT 1953.230 30.840 1953.550 30.900 ;
        RECT 1347.410 30.700 1953.550 30.840 ;
        RECT 1347.410 30.640 1347.730 30.700 ;
        RECT 1953.230 30.640 1953.550 30.700 ;
      LAYER via ;
        RECT 1347.900 1684.060 1348.160 1684.320 ;
        RECT 1350.660 1684.060 1350.920 1684.320 ;
        RECT 1347.900 1634.760 1348.160 1635.020 ;
        RECT 1347.440 1633.740 1347.700 1634.000 ;
        RECT 1347.440 30.640 1347.700 30.900 ;
        RECT 1953.260 30.640 1953.520 30.900 ;
      LAYER met2 ;
        RECT 1350.560 1700.340 1350.840 1704.000 ;
        RECT 1350.560 1700.000 1350.860 1700.340 ;
        RECT 1350.720 1684.350 1350.860 1700.000 ;
        RECT 1347.900 1684.030 1348.160 1684.350 ;
        RECT 1350.660 1684.030 1350.920 1684.350 ;
        RECT 1347.960 1635.050 1348.100 1684.030 ;
        RECT 1347.900 1634.730 1348.160 1635.050 ;
        RECT 1347.440 1633.710 1347.700 1634.030 ;
        RECT 1347.500 30.930 1347.640 1633.710 ;
        RECT 1347.440 30.610 1347.700 30.930 ;
        RECT 1953.260 30.610 1953.520 30.930 ;
        RECT 1953.320 2.400 1953.460 30.610 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1352.470 1654.000 1352.790 1654.060 ;
        RECT 1966.570 1654.000 1966.890 1654.060 ;
        RECT 1352.470 1653.860 1966.890 1654.000 ;
        RECT 1352.470 1653.800 1352.790 1653.860 ;
        RECT 1966.570 1653.800 1966.890 1653.860 ;
      LAYER via ;
        RECT 1352.500 1653.800 1352.760 1654.060 ;
        RECT 1966.600 1653.800 1966.860 1654.060 ;
      LAYER met2 ;
        RECT 1352.400 1700.340 1352.680 1704.000 ;
        RECT 1352.400 1700.000 1352.700 1700.340 ;
        RECT 1352.560 1654.090 1352.700 1700.000 ;
        RECT 1352.500 1653.770 1352.760 1654.090 ;
        RECT 1966.600 1653.770 1966.860 1654.090 ;
        RECT 1966.660 17.410 1966.800 1653.770 ;
        RECT 1966.660 17.270 1971.400 17.410 ;
        RECT 1971.260 2.400 1971.400 17.270 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1386.585 1676.625 1386.755 1690.735 ;
      LAYER mcon ;
        RECT 1386.585 1690.565 1386.755 1690.735 ;
      LAYER met1 ;
        RECT 1354.310 1690.720 1354.630 1690.780 ;
        RECT 1386.525 1690.720 1386.815 1690.765 ;
        RECT 1354.310 1690.580 1386.815 1690.720 ;
        RECT 1354.310 1690.520 1354.630 1690.580 ;
        RECT 1386.525 1690.535 1386.815 1690.580 ;
        RECT 1386.525 1676.780 1386.815 1676.825 ;
        RECT 1401.690 1676.780 1402.010 1676.840 ;
        RECT 1386.525 1676.640 1402.010 1676.780 ;
        RECT 1386.525 1676.595 1386.815 1676.640 ;
        RECT 1401.690 1676.580 1402.010 1676.640 ;
        RECT 1401.690 1646.520 1402.010 1646.580 ;
        RECT 1987.270 1646.520 1987.590 1646.580 ;
        RECT 1401.690 1646.380 1987.590 1646.520 ;
        RECT 1401.690 1646.320 1402.010 1646.380 ;
        RECT 1987.270 1646.320 1987.590 1646.380 ;
      LAYER via ;
        RECT 1354.340 1690.520 1354.600 1690.780 ;
        RECT 1401.720 1676.580 1401.980 1676.840 ;
        RECT 1401.720 1646.320 1401.980 1646.580 ;
        RECT 1987.300 1646.320 1987.560 1646.580 ;
      LAYER met2 ;
        RECT 1354.240 1700.340 1354.520 1704.000 ;
        RECT 1354.240 1700.000 1354.540 1700.340 ;
        RECT 1354.400 1690.810 1354.540 1700.000 ;
        RECT 1354.340 1690.490 1354.600 1690.810 ;
        RECT 1401.720 1676.550 1401.980 1676.870 ;
        RECT 1401.780 1646.610 1401.920 1676.550 ;
        RECT 1401.720 1646.290 1401.980 1646.610 ;
        RECT 1987.300 1646.290 1987.560 1646.610 ;
        RECT 1987.360 17.410 1987.500 1646.290 ;
        RECT 1987.360 17.270 1989.340 17.410 ;
        RECT 1989.200 2.400 1989.340 17.270 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1356.150 1667.260 1356.470 1667.320 ;
        RECT 2001.530 1667.260 2001.850 1667.320 ;
        RECT 1356.150 1667.120 2001.850 1667.260 ;
        RECT 1356.150 1667.060 1356.470 1667.120 ;
        RECT 2001.530 1667.060 2001.850 1667.120 ;
      LAYER via ;
        RECT 1356.180 1667.060 1356.440 1667.320 ;
        RECT 2001.560 1667.060 2001.820 1667.320 ;
      LAYER met2 ;
        RECT 1356.080 1700.340 1356.360 1704.000 ;
        RECT 1356.080 1700.000 1356.380 1700.340 ;
        RECT 1356.240 1667.350 1356.380 1700.000 ;
        RECT 1356.180 1667.030 1356.440 1667.350 ;
        RECT 2001.560 1667.030 2001.820 1667.350 ;
        RECT 2001.620 17.410 2001.760 1667.030 ;
        RECT 2001.620 17.270 2006.820 17.410 ;
        RECT 2006.680 2.400 2006.820 17.270 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1357.990 1660.460 1358.310 1660.520 ;
        RECT 2021.770 1660.460 2022.090 1660.520 ;
        RECT 1357.990 1660.320 2022.090 1660.460 ;
        RECT 1357.990 1660.260 1358.310 1660.320 ;
        RECT 2021.770 1660.260 2022.090 1660.320 ;
      LAYER via ;
        RECT 1358.020 1660.260 1358.280 1660.520 ;
        RECT 2021.800 1660.260 2022.060 1660.520 ;
      LAYER met2 ;
        RECT 1357.920 1700.340 1358.200 1704.000 ;
        RECT 1357.920 1700.000 1358.220 1700.340 ;
        RECT 1358.080 1660.550 1358.220 1700.000 ;
        RECT 1358.020 1660.230 1358.280 1660.550 ;
        RECT 2021.800 1660.230 2022.060 1660.550 ;
        RECT 2021.860 17.410 2022.000 1660.230 ;
        RECT 2021.860 17.270 2024.760 17.410 ;
        RECT 2024.620 2.400 2024.760 17.270 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1365.885 1688.865 1366.055 1690.055 ;
        RECT 1379.685 1687.505 1379.855 1689.035 ;
      LAYER mcon ;
        RECT 1365.885 1689.885 1366.055 1690.055 ;
        RECT 1379.685 1688.865 1379.855 1689.035 ;
      LAYER met1 ;
        RECT 1359.830 1690.380 1360.150 1690.440 ;
        RECT 1359.830 1690.240 1366.040 1690.380 ;
        RECT 1359.830 1690.180 1360.150 1690.240 ;
        RECT 1365.900 1690.085 1366.040 1690.240 ;
        RECT 1365.825 1689.855 1366.115 1690.085 ;
        RECT 1365.825 1689.020 1366.115 1689.065 ;
        RECT 1379.625 1689.020 1379.915 1689.065 ;
        RECT 1365.825 1688.880 1379.915 1689.020 ;
        RECT 1365.825 1688.835 1366.115 1688.880 ;
        RECT 1379.625 1688.835 1379.915 1688.880 ;
        RECT 1379.625 1687.660 1379.915 1687.705 ;
        RECT 1415.030 1687.660 1415.350 1687.720 ;
        RECT 1379.625 1687.520 1415.350 1687.660 ;
        RECT 1379.625 1687.475 1379.915 1687.520 ;
        RECT 1415.030 1687.460 1415.350 1687.520 ;
        RECT 1414.570 1676.780 1414.890 1676.840 ;
        RECT 1416.410 1676.780 1416.730 1676.840 ;
        RECT 1414.570 1676.640 1416.730 1676.780 ;
        RECT 1414.570 1676.580 1414.890 1676.640 ;
        RECT 1416.410 1676.580 1416.730 1676.640 ;
        RECT 1416.410 1639.720 1416.730 1639.780 ;
        RECT 2042.470 1639.720 2042.790 1639.780 ;
        RECT 1416.410 1639.580 2042.790 1639.720 ;
        RECT 1416.410 1639.520 1416.730 1639.580 ;
        RECT 2042.470 1639.520 2042.790 1639.580 ;
      LAYER via ;
        RECT 1359.860 1690.180 1360.120 1690.440 ;
        RECT 1415.060 1687.460 1415.320 1687.720 ;
        RECT 1414.600 1676.580 1414.860 1676.840 ;
        RECT 1416.440 1676.580 1416.700 1676.840 ;
        RECT 1416.440 1639.520 1416.700 1639.780 ;
        RECT 2042.500 1639.520 2042.760 1639.780 ;
      LAYER met2 ;
        RECT 1359.760 1700.340 1360.040 1704.000 ;
        RECT 1359.760 1700.000 1360.060 1700.340 ;
        RECT 1359.920 1690.470 1360.060 1700.000 ;
        RECT 1359.860 1690.150 1360.120 1690.470 ;
        RECT 1415.060 1687.430 1415.320 1687.750 ;
        RECT 1415.120 1683.410 1415.260 1687.430 ;
        RECT 1414.660 1683.270 1415.260 1683.410 ;
        RECT 1414.660 1676.870 1414.800 1683.270 ;
        RECT 1414.600 1676.550 1414.860 1676.870 ;
        RECT 1416.440 1676.550 1416.700 1676.870 ;
        RECT 1416.500 1639.810 1416.640 1676.550 ;
        RECT 1416.440 1639.490 1416.700 1639.810 ;
        RECT 2042.500 1639.490 2042.760 1639.810 ;
        RECT 2042.560 2.400 2042.700 1639.490 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1221.830 1663.180 1222.150 1663.240 ;
        RECT 1227.350 1663.180 1227.670 1663.240 ;
        RECT 1221.830 1663.040 1227.670 1663.180 ;
        RECT 1221.830 1662.980 1222.150 1663.040 ;
        RECT 1227.350 1662.980 1227.670 1663.040 ;
        RECT 758.610 1653.660 758.930 1653.720 ;
        RECT 1221.830 1653.660 1222.150 1653.720 ;
        RECT 758.610 1653.520 1222.150 1653.660 ;
        RECT 758.610 1653.460 758.930 1653.520 ;
        RECT 1221.830 1653.460 1222.150 1653.520 ;
      LAYER via ;
        RECT 1221.860 1662.980 1222.120 1663.240 ;
        RECT 1227.380 1662.980 1227.640 1663.240 ;
        RECT 758.640 1653.460 758.900 1653.720 ;
        RECT 1221.860 1653.460 1222.120 1653.720 ;
      LAYER met2 ;
        RECT 1227.280 1700.340 1227.560 1704.000 ;
        RECT 1227.280 1700.000 1227.580 1700.340 ;
        RECT 1227.440 1663.270 1227.580 1700.000 ;
        RECT 1221.860 1662.950 1222.120 1663.270 ;
        RECT 1227.380 1662.950 1227.640 1663.270 ;
        RECT 1221.920 1653.750 1222.060 1662.950 ;
        RECT 758.640 1653.430 758.900 1653.750 ;
        RECT 1221.860 1653.430 1222.120 1653.750 ;
        RECT 758.700 17.410 758.840 1653.430 ;
        RECT 757.780 17.270 758.840 17.410 ;
        RECT 757.780 2.400 757.920 17.270 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1361.670 1683.920 1361.990 1683.980 ;
        RECT 1363.050 1683.920 1363.370 1683.980 ;
        RECT 1361.670 1683.780 1363.370 1683.920 ;
        RECT 1361.670 1683.720 1361.990 1683.780 ;
        RECT 1363.050 1683.720 1363.370 1683.780 ;
        RECT 1363.050 1653.660 1363.370 1653.720 ;
        RECT 2056.270 1653.660 2056.590 1653.720 ;
        RECT 1363.050 1653.520 2056.590 1653.660 ;
        RECT 1363.050 1653.460 1363.370 1653.520 ;
        RECT 2056.270 1653.460 2056.590 1653.520 ;
      LAYER via ;
        RECT 1361.700 1683.720 1361.960 1683.980 ;
        RECT 1363.080 1683.720 1363.340 1683.980 ;
        RECT 1363.080 1653.460 1363.340 1653.720 ;
        RECT 2056.300 1653.460 2056.560 1653.720 ;
      LAYER met2 ;
        RECT 1361.600 1700.340 1361.880 1704.000 ;
        RECT 1361.600 1700.000 1361.900 1700.340 ;
        RECT 1361.760 1684.010 1361.900 1700.000 ;
        RECT 1361.700 1683.690 1361.960 1684.010 ;
        RECT 1363.080 1683.690 1363.340 1684.010 ;
        RECT 1363.140 1653.750 1363.280 1683.690 ;
        RECT 1363.080 1653.430 1363.340 1653.750 ;
        RECT 2056.300 1653.430 2056.560 1653.750 ;
        RECT 2056.360 17.410 2056.500 1653.430 ;
        RECT 2056.360 17.270 2060.640 17.410 ;
        RECT 2060.500 2.400 2060.640 17.270 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1545.745 1632.765 1547.295 1632.935 ;
      LAYER mcon ;
        RECT 1547.125 1632.765 1547.295 1632.935 ;
      LAYER met1 ;
        RECT 1363.510 1683.920 1363.830 1683.980 ;
        RECT 1363.510 1683.780 1364.200 1683.920 ;
        RECT 1363.510 1683.720 1363.830 1683.780 ;
        RECT 1364.060 1683.240 1364.200 1683.780 ;
        RECT 1365.350 1683.240 1365.670 1683.300 ;
        RECT 1364.060 1683.100 1365.670 1683.240 ;
        RECT 1365.350 1683.040 1365.670 1683.100 ;
        RECT 1365.350 1632.920 1365.670 1632.980 ;
        RECT 1545.685 1632.920 1545.975 1632.965 ;
        RECT 1365.350 1632.780 1545.975 1632.920 ;
        RECT 1365.350 1632.720 1365.670 1632.780 ;
        RECT 1545.685 1632.735 1545.975 1632.780 ;
        RECT 1547.065 1632.920 1547.355 1632.965 ;
        RECT 2076.970 1632.920 2077.290 1632.980 ;
        RECT 1547.065 1632.780 2077.290 1632.920 ;
        RECT 1547.065 1632.735 1547.355 1632.780 ;
        RECT 2076.970 1632.720 2077.290 1632.780 ;
      LAYER via ;
        RECT 1363.540 1683.720 1363.800 1683.980 ;
        RECT 1365.380 1683.040 1365.640 1683.300 ;
        RECT 1365.380 1632.720 1365.640 1632.980 ;
        RECT 2077.000 1632.720 2077.260 1632.980 ;
      LAYER met2 ;
        RECT 1363.440 1700.340 1363.720 1704.000 ;
        RECT 1363.440 1700.000 1363.740 1700.340 ;
        RECT 1363.600 1684.010 1363.740 1700.000 ;
        RECT 1363.540 1683.690 1363.800 1684.010 ;
        RECT 1365.380 1683.010 1365.640 1683.330 ;
        RECT 1365.440 1633.010 1365.580 1683.010 ;
        RECT 1365.380 1632.690 1365.640 1633.010 ;
        RECT 2077.000 1632.690 2077.260 1633.010 ;
        RECT 2077.060 17.410 2077.200 1632.690 ;
        RECT 2077.060 17.270 2078.580 17.410 ;
        RECT 2078.440 2.400 2078.580 17.270 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1364.430 1683.920 1364.750 1683.980 ;
        RECT 1365.350 1683.920 1365.670 1683.980 ;
        RECT 1364.430 1683.780 1365.670 1683.920 ;
        RECT 1364.430 1683.720 1364.750 1683.780 ;
        RECT 1365.350 1683.720 1365.670 1683.780 ;
        RECT 1364.430 1625.440 1364.750 1625.500 ;
        RECT 2090.770 1625.440 2091.090 1625.500 ;
        RECT 1364.430 1625.300 2091.090 1625.440 ;
        RECT 1364.430 1625.240 1364.750 1625.300 ;
        RECT 2090.770 1625.240 2091.090 1625.300 ;
      LAYER via ;
        RECT 1364.460 1683.720 1364.720 1683.980 ;
        RECT 1365.380 1683.720 1365.640 1683.980 ;
        RECT 1364.460 1625.240 1364.720 1625.500 ;
        RECT 2090.800 1625.240 2091.060 1625.500 ;
      LAYER met2 ;
        RECT 1365.280 1700.340 1365.560 1704.000 ;
        RECT 1365.280 1700.000 1365.580 1700.340 ;
        RECT 1365.440 1684.010 1365.580 1700.000 ;
        RECT 1364.460 1683.690 1364.720 1684.010 ;
        RECT 1365.380 1683.690 1365.640 1684.010 ;
        RECT 1364.520 1625.530 1364.660 1683.690 ;
        RECT 1364.460 1625.210 1364.720 1625.530 ;
        RECT 2090.800 1625.210 2091.060 1625.530 ;
        RECT 2090.860 17.410 2091.000 1625.210 ;
        RECT 2090.860 17.270 2096.060 17.410 ;
        RECT 2095.920 2.400 2096.060 17.270 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1366.270 1686.980 1366.590 1687.040 ;
        RECT 1367.190 1686.980 1367.510 1687.040 ;
        RECT 1366.270 1686.840 1367.510 1686.980 ;
        RECT 1366.270 1686.780 1366.590 1686.840 ;
        RECT 1367.190 1686.780 1367.510 1686.840 ;
        RECT 1366.270 1674.060 1366.590 1674.120 ;
        RECT 2111.470 1674.060 2111.790 1674.120 ;
        RECT 1366.270 1673.920 2111.790 1674.060 ;
        RECT 1366.270 1673.860 1366.590 1673.920 ;
        RECT 2111.470 1673.860 2111.790 1673.920 ;
      LAYER via ;
        RECT 1366.300 1686.780 1366.560 1687.040 ;
        RECT 1367.220 1686.780 1367.480 1687.040 ;
        RECT 1366.300 1673.860 1366.560 1674.120 ;
        RECT 2111.500 1673.860 2111.760 1674.120 ;
      LAYER met2 ;
        RECT 1367.120 1700.340 1367.400 1704.000 ;
        RECT 1367.120 1700.000 1367.420 1700.340 ;
        RECT 1367.280 1687.070 1367.420 1700.000 ;
        RECT 1366.300 1686.750 1366.560 1687.070 ;
        RECT 1367.220 1686.750 1367.480 1687.070 ;
        RECT 1366.360 1674.150 1366.500 1686.750 ;
        RECT 1366.300 1673.830 1366.560 1674.150 ;
        RECT 2111.500 1673.830 2111.760 1674.150 ;
        RECT 2111.560 17.410 2111.700 1673.830 ;
        RECT 2111.560 17.270 2114.000 17.410 ;
        RECT 2113.860 2.400 2114.000 17.270 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1366.730 1684.600 1367.050 1684.660 ;
        RECT 1369.030 1684.600 1369.350 1684.660 ;
        RECT 1366.730 1684.460 1369.350 1684.600 ;
        RECT 1366.730 1684.400 1367.050 1684.460 ;
        RECT 1369.030 1684.400 1369.350 1684.460 ;
        RECT 1366.730 1646.180 1367.050 1646.240 ;
        RECT 2125.730 1646.180 2126.050 1646.240 ;
        RECT 1366.730 1646.040 2126.050 1646.180 ;
        RECT 1366.730 1645.980 1367.050 1646.040 ;
        RECT 2125.730 1645.980 2126.050 1646.040 ;
        RECT 2125.730 14.520 2126.050 14.580 ;
        RECT 2131.710 14.520 2132.030 14.580 ;
        RECT 2125.730 14.380 2132.030 14.520 ;
        RECT 2125.730 14.320 2126.050 14.380 ;
        RECT 2131.710 14.320 2132.030 14.380 ;
      LAYER via ;
        RECT 1366.760 1684.400 1367.020 1684.660 ;
        RECT 1369.060 1684.400 1369.320 1684.660 ;
        RECT 1366.760 1645.980 1367.020 1646.240 ;
        RECT 2125.760 1645.980 2126.020 1646.240 ;
        RECT 2125.760 14.320 2126.020 14.580 ;
        RECT 2131.740 14.320 2132.000 14.580 ;
      LAYER met2 ;
        RECT 1368.960 1700.340 1369.240 1704.000 ;
        RECT 1368.960 1700.000 1369.260 1700.340 ;
        RECT 1369.120 1684.690 1369.260 1700.000 ;
        RECT 1366.760 1684.370 1367.020 1684.690 ;
        RECT 1369.060 1684.370 1369.320 1684.690 ;
        RECT 1366.820 1646.270 1366.960 1684.370 ;
        RECT 1366.760 1645.950 1367.020 1646.270 ;
        RECT 2125.760 1645.950 2126.020 1646.270 ;
        RECT 2125.820 14.610 2125.960 1645.950 ;
        RECT 2125.760 14.290 2126.020 14.610 ;
        RECT 2131.740 14.290 2132.000 14.610 ;
        RECT 2131.800 2.400 2131.940 14.290 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1368.110 1684.260 1368.430 1684.320 ;
        RECT 1370.870 1684.260 1371.190 1684.320 ;
        RECT 1368.110 1684.120 1371.190 1684.260 ;
        RECT 1368.110 1684.060 1368.430 1684.120 ;
        RECT 1370.870 1684.060 1371.190 1684.120 ;
        RECT 1368.110 1639.380 1368.430 1639.440 ;
        RECT 2145.970 1639.380 2146.290 1639.440 ;
        RECT 1368.110 1639.240 2146.290 1639.380 ;
        RECT 1368.110 1639.180 1368.430 1639.240 ;
        RECT 2145.970 1639.180 2146.290 1639.240 ;
      LAYER via ;
        RECT 1368.140 1684.060 1368.400 1684.320 ;
        RECT 1370.900 1684.060 1371.160 1684.320 ;
        RECT 1368.140 1639.180 1368.400 1639.440 ;
        RECT 2146.000 1639.180 2146.260 1639.440 ;
      LAYER met2 ;
        RECT 1370.800 1700.340 1371.080 1704.000 ;
        RECT 1370.800 1700.000 1371.100 1700.340 ;
        RECT 1370.960 1684.350 1371.100 1700.000 ;
        RECT 1368.140 1684.030 1368.400 1684.350 ;
        RECT 1370.900 1684.030 1371.160 1684.350 ;
        RECT 1368.200 1639.470 1368.340 1684.030 ;
        RECT 1368.140 1639.150 1368.400 1639.470 ;
        RECT 2146.000 1639.150 2146.260 1639.470 ;
        RECT 2146.060 17.410 2146.200 1639.150 ;
        RECT 2146.060 17.270 2149.880 17.410 ;
        RECT 2149.740 2.400 2149.880 17.270 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1372.710 1597.900 1373.030 1597.960 ;
        RECT 2167.130 1597.900 2167.450 1597.960 ;
        RECT 1372.710 1597.760 2167.450 1597.900 ;
        RECT 1372.710 1597.700 1373.030 1597.760 ;
        RECT 2167.130 1597.700 2167.450 1597.760 ;
      LAYER via ;
        RECT 1372.740 1597.700 1373.000 1597.960 ;
        RECT 2167.160 1597.700 2167.420 1597.960 ;
      LAYER met2 ;
        RECT 1372.640 1700.340 1372.920 1704.000 ;
        RECT 1372.640 1700.000 1372.940 1700.340 ;
        RECT 1372.800 1597.990 1372.940 1700.000 ;
        RECT 1372.740 1597.670 1373.000 1597.990 ;
        RECT 2167.160 1597.670 2167.420 1597.990 ;
        RECT 2167.220 17.410 2167.360 1597.670 ;
        RECT 2167.220 17.270 2167.820 17.410 ;
        RECT 2167.680 2.400 2167.820 17.270 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1374.550 1685.280 1374.870 1685.340 ;
        RECT 1374.550 1685.140 1387.200 1685.280 ;
        RECT 1374.550 1685.080 1374.870 1685.140 ;
        RECT 1387.060 1683.920 1387.200 1685.140 ;
        RECT 1387.060 1683.780 1387.660 1683.920 ;
        RECT 1387.520 1683.580 1387.660 1683.780 ;
        RECT 1393.410 1683.580 1393.730 1683.640 ;
        RECT 1387.520 1683.440 1393.730 1683.580 ;
        RECT 1393.410 1683.380 1393.730 1683.440 ;
        RECT 1393.870 1676.100 1394.190 1676.160 ;
        RECT 1395.710 1676.100 1396.030 1676.160 ;
        RECT 1393.870 1675.960 1396.030 1676.100 ;
        RECT 1393.870 1675.900 1394.190 1675.960 ;
        RECT 1395.710 1675.900 1396.030 1675.960 ;
        RECT 1395.710 1618.980 1396.030 1619.040 ;
        RECT 2180.470 1618.980 2180.790 1619.040 ;
        RECT 1395.710 1618.840 2180.790 1618.980 ;
        RECT 1395.710 1618.780 1396.030 1618.840 ;
        RECT 2180.470 1618.780 2180.790 1618.840 ;
      LAYER via ;
        RECT 1374.580 1685.080 1374.840 1685.340 ;
        RECT 1393.440 1683.380 1393.700 1683.640 ;
        RECT 1393.900 1675.900 1394.160 1676.160 ;
        RECT 1395.740 1675.900 1396.000 1676.160 ;
        RECT 1395.740 1618.780 1396.000 1619.040 ;
        RECT 2180.500 1618.780 2180.760 1619.040 ;
      LAYER met2 ;
        RECT 1374.480 1700.340 1374.760 1704.000 ;
        RECT 1374.480 1700.000 1374.780 1700.340 ;
        RECT 1374.640 1685.370 1374.780 1700.000 ;
        RECT 1374.580 1685.050 1374.840 1685.370 ;
        RECT 1393.440 1683.350 1393.700 1683.670 ;
        RECT 1393.500 1682.050 1393.640 1683.350 ;
        RECT 1393.500 1681.910 1394.100 1682.050 ;
        RECT 1393.960 1676.190 1394.100 1681.910 ;
        RECT 1393.900 1675.870 1394.160 1676.190 ;
        RECT 1395.740 1675.870 1396.000 1676.190 ;
        RECT 1395.800 1619.070 1395.940 1675.870 ;
        RECT 1395.740 1618.750 1396.000 1619.070 ;
        RECT 2180.500 1618.750 2180.760 1619.070 ;
        RECT 2180.560 17.410 2180.700 1618.750 ;
        RECT 2180.560 17.270 2185.300 17.410 ;
        RECT 2185.160 2.400 2185.300 17.270 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1376.390 1684.940 1376.710 1685.000 ;
        RECT 1377.770 1684.940 1378.090 1685.000 ;
        RECT 1376.390 1684.800 1378.090 1684.940 ;
        RECT 1376.390 1684.740 1376.710 1684.800 ;
        RECT 1377.770 1684.740 1378.090 1684.800 ;
        RECT 1377.770 1666.920 1378.090 1666.980 ;
        RECT 2201.170 1666.920 2201.490 1666.980 ;
        RECT 1377.770 1666.780 2201.490 1666.920 ;
        RECT 1377.770 1666.720 1378.090 1666.780 ;
        RECT 2201.170 1666.720 2201.490 1666.780 ;
      LAYER via ;
        RECT 1376.420 1684.740 1376.680 1685.000 ;
        RECT 1377.800 1684.740 1378.060 1685.000 ;
        RECT 1377.800 1666.720 1378.060 1666.980 ;
        RECT 2201.200 1666.720 2201.460 1666.980 ;
      LAYER met2 ;
        RECT 1376.320 1700.340 1376.600 1704.000 ;
        RECT 1376.320 1700.000 1376.620 1700.340 ;
        RECT 1376.480 1685.030 1376.620 1700.000 ;
        RECT 1376.420 1684.710 1376.680 1685.030 ;
        RECT 1377.800 1684.710 1378.060 1685.030 ;
        RECT 1377.860 1667.010 1378.000 1684.710 ;
        RECT 1377.800 1666.690 1378.060 1667.010 ;
        RECT 2201.200 1666.690 2201.460 1667.010 ;
        RECT 2201.260 17.410 2201.400 1666.690 ;
        RECT 2201.260 17.270 2203.240 17.410 ;
        RECT 2203.100 2.400 2203.240 17.270 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1378.230 1681.200 1378.550 1681.260 ;
        RECT 2215.430 1681.200 2215.750 1681.260 ;
        RECT 1378.230 1681.060 2215.750 1681.200 ;
        RECT 1378.230 1681.000 1378.550 1681.060 ;
        RECT 2215.430 1681.000 2215.750 1681.060 ;
      LAYER via ;
        RECT 1378.260 1681.000 1378.520 1681.260 ;
        RECT 2215.460 1681.000 2215.720 1681.260 ;
      LAYER met2 ;
        RECT 1378.160 1700.340 1378.440 1704.000 ;
        RECT 1378.160 1700.000 1378.460 1700.340 ;
        RECT 1378.320 1681.290 1378.460 1700.000 ;
        RECT 1378.260 1680.970 1378.520 1681.290 ;
        RECT 2215.460 1680.970 2215.720 1681.290 ;
        RECT 2215.520 17.410 2215.660 1680.970 ;
        RECT 2215.520 17.270 2221.180 17.410 ;
        RECT 2221.040 2.400 2221.180 17.270 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1221.370 1683.920 1221.690 1683.980 ;
        RECT 1229.190 1683.920 1229.510 1683.980 ;
        RECT 1221.370 1683.780 1229.510 1683.920 ;
        RECT 1221.370 1683.720 1221.690 1683.780 ;
        RECT 1229.190 1683.720 1229.510 1683.780 ;
        RECT 779.310 1646.180 779.630 1646.240 ;
        RECT 1221.370 1646.180 1221.690 1646.240 ;
        RECT 779.310 1646.040 1221.690 1646.180 ;
        RECT 779.310 1645.980 779.630 1646.040 ;
        RECT 1221.370 1645.980 1221.690 1646.040 ;
      LAYER via ;
        RECT 1221.400 1683.720 1221.660 1683.980 ;
        RECT 1229.220 1683.720 1229.480 1683.980 ;
        RECT 779.340 1645.980 779.600 1646.240 ;
        RECT 1221.400 1645.980 1221.660 1646.240 ;
      LAYER met2 ;
        RECT 1229.120 1700.340 1229.400 1704.000 ;
        RECT 1229.120 1700.000 1229.420 1700.340 ;
        RECT 1229.280 1684.010 1229.420 1700.000 ;
        RECT 1221.400 1683.690 1221.660 1684.010 ;
        RECT 1229.220 1683.690 1229.480 1684.010 ;
        RECT 1221.460 1646.270 1221.600 1683.690 ;
        RECT 779.340 1645.950 779.600 1646.270 ;
        RECT 1221.400 1645.950 1221.660 1646.270 ;
        RECT 779.400 18.090 779.540 1645.950 ;
        RECT 775.720 17.950 779.540 18.090 ;
        RECT 775.720 2.400 775.860 17.950 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1402.685 1676.625 1402.855 1688.695 ;
      LAYER mcon ;
        RECT 1402.685 1688.525 1402.855 1688.695 ;
      LAYER met1 ;
        RECT 1380.070 1689.020 1380.390 1689.080 ;
        RECT 1380.070 1688.880 1400.080 1689.020 ;
        RECT 1380.070 1688.820 1380.390 1688.880 ;
        RECT 1399.940 1688.680 1400.080 1688.880 ;
        RECT 1402.625 1688.680 1402.915 1688.725 ;
        RECT 1399.940 1688.540 1402.915 1688.680 ;
        RECT 1402.625 1688.495 1402.915 1688.540 ;
        RECT 1402.610 1676.780 1402.930 1676.840 ;
        RECT 1402.415 1676.640 1402.930 1676.780 ;
        RECT 1402.610 1676.580 1402.930 1676.640 ;
        RECT 1402.610 1590.760 1402.930 1590.820 ;
        RECT 2235.670 1590.760 2235.990 1590.820 ;
        RECT 1402.610 1590.620 2235.990 1590.760 ;
        RECT 1402.610 1590.560 1402.930 1590.620 ;
        RECT 2235.670 1590.560 2235.990 1590.620 ;
      LAYER via ;
        RECT 1380.100 1688.820 1380.360 1689.080 ;
        RECT 1402.640 1676.580 1402.900 1676.840 ;
        RECT 1402.640 1590.560 1402.900 1590.820 ;
        RECT 2235.700 1590.560 2235.960 1590.820 ;
      LAYER met2 ;
        RECT 1380.000 1700.340 1380.280 1704.000 ;
        RECT 1380.000 1700.000 1380.300 1700.340 ;
        RECT 1380.160 1689.110 1380.300 1700.000 ;
        RECT 1380.100 1688.790 1380.360 1689.110 ;
        RECT 1402.640 1676.550 1402.900 1676.870 ;
        RECT 1402.700 1590.850 1402.840 1676.550 ;
        RECT 1402.640 1590.530 1402.900 1590.850 ;
        RECT 2235.700 1590.530 2235.960 1590.850 ;
        RECT 2235.760 17.410 2235.900 1590.530 ;
        RECT 2235.760 17.270 2239.120 17.410 ;
        RECT 2238.980 2.400 2239.120 17.270 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1381.910 1678.480 1382.230 1678.540 ;
        RECT 1386.050 1678.480 1386.370 1678.540 ;
        RECT 1381.910 1678.340 1386.370 1678.480 ;
        RECT 1381.910 1678.280 1382.230 1678.340 ;
        RECT 1386.050 1678.280 1386.370 1678.340 ;
        RECT 1386.050 1653.320 1386.370 1653.380 ;
        RECT 2256.370 1653.320 2256.690 1653.380 ;
        RECT 1386.050 1653.180 2256.690 1653.320 ;
        RECT 1386.050 1653.120 1386.370 1653.180 ;
        RECT 2256.370 1653.120 2256.690 1653.180 ;
      LAYER via ;
        RECT 1381.940 1678.280 1382.200 1678.540 ;
        RECT 1386.080 1678.280 1386.340 1678.540 ;
        RECT 1386.080 1653.120 1386.340 1653.380 ;
        RECT 2256.400 1653.120 2256.660 1653.380 ;
      LAYER met2 ;
        RECT 1381.840 1700.340 1382.120 1704.000 ;
        RECT 1381.840 1700.000 1382.140 1700.340 ;
        RECT 1382.000 1678.570 1382.140 1700.000 ;
        RECT 1381.940 1678.250 1382.200 1678.570 ;
        RECT 1386.080 1678.250 1386.340 1678.570 ;
        RECT 1386.140 1653.410 1386.280 1678.250 ;
        RECT 1386.080 1653.090 1386.340 1653.410 ;
        RECT 2256.400 1653.090 2256.660 1653.410 ;
        RECT 2256.460 2.400 2256.600 1653.090 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1383.750 1611.840 1384.070 1611.900 ;
        RECT 2270.170 1611.840 2270.490 1611.900 ;
        RECT 1383.750 1611.700 2270.490 1611.840 ;
        RECT 1383.750 1611.640 1384.070 1611.700 ;
        RECT 2270.170 1611.640 2270.490 1611.700 ;
      LAYER via ;
        RECT 1383.780 1611.640 1384.040 1611.900 ;
        RECT 2270.200 1611.640 2270.460 1611.900 ;
      LAYER met2 ;
        RECT 1383.680 1700.340 1383.960 1704.000 ;
        RECT 1383.680 1700.000 1383.980 1700.340 ;
        RECT 1383.840 1611.930 1383.980 1700.000 ;
        RECT 1383.780 1611.610 1384.040 1611.930 ;
        RECT 2270.200 1611.610 2270.460 1611.930 ;
        RECT 2270.260 17.410 2270.400 1611.610 ;
        RECT 2270.260 17.270 2274.540 17.410 ;
        RECT 2274.400 2.400 2274.540 17.270 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1380.990 1684.260 1381.310 1684.320 ;
        RECT 1385.590 1684.260 1385.910 1684.320 ;
        RECT 1380.990 1684.120 1385.910 1684.260 ;
        RECT 1380.990 1684.060 1381.310 1684.120 ;
        RECT 1385.590 1684.060 1385.910 1684.120 ;
        RECT 1381.450 1583.960 1381.770 1584.020 ;
        RECT 2290.870 1583.960 2291.190 1584.020 ;
        RECT 1381.450 1583.820 2291.190 1583.960 ;
        RECT 1381.450 1583.760 1381.770 1583.820 ;
        RECT 2290.870 1583.760 2291.190 1583.820 ;
      LAYER via ;
        RECT 1381.020 1684.060 1381.280 1684.320 ;
        RECT 1385.620 1684.060 1385.880 1684.320 ;
        RECT 1381.480 1583.760 1381.740 1584.020 ;
        RECT 2290.900 1583.760 2291.160 1584.020 ;
      LAYER met2 ;
        RECT 1385.520 1700.340 1385.800 1704.000 ;
        RECT 1385.520 1700.000 1385.820 1700.340 ;
        RECT 1385.680 1684.350 1385.820 1700.000 ;
        RECT 1381.020 1684.030 1381.280 1684.350 ;
        RECT 1385.620 1684.030 1385.880 1684.350 ;
        RECT 1381.080 1666.410 1381.220 1684.030 ;
        RECT 1381.080 1666.270 1381.680 1666.410 ;
        RECT 1381.540 1584.050 1381.680 1666.270 ;
        RECT 1381.480 1583.730 1381.740 1584.050 ;
        RECT 2290.900 1583.730 2291.160 1584.050 ;
        RECT 2290.960 17.410 2291.100 1583.730 ;
        RECT 2290.960 17.270 2292.480 17.410 ;
        RECT 2292.340 2.400 2292.480 17.270 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1404.985 1675.945 1405.155 1689.375 ;
      LAYER mcon ;
        RECT 1404.985 1689.205 1405.155 1689.375 ;
      LAYER met1 ;
        RECT 1387.430 1689.360 1387.750 1689.420 ;
        RECT 1404.925 1689.360 1405.215 1689.405 ;
        RECT 1387.430 1689.220 1405.215 1689.360 ;
        RECT 1387.430 1689.160 1387.750 1689.220 ;
        RECT 1404.925 1689.175 1405.215 1689.220 ;
        RECT 1404.925 1676.100 1405.215 1676.145 ;
        RECT 1417.330 1676.100 1417.650 1676.160 ;
        RECT 1404.925 1675.960 1417.650 1676.100 ;
        RECT 1404.925 1675.915 1405.215 1675.960 ;
        RECT 1417.330 1675.900 1417.650 1675.960 ;
        RECT 1417.330 1576.820 1417.650 1576.880 ;
        RECT 2304.670 1576.820 2304.990 1576.880 ;
        RECT 1417.330 1576.680 2304.990 1576.820 ;
        RECT 1417.330 1576.620 1417.650 1576.680 ;
        RECT 2304.670 1576.620 2304.990 1576.680 ;
      LAYER via ;
        RECT 1387.460 1689.160 1387.720 1689.420 ;
        RECT 1417.360 1675.900 1417.620 1676.160 ;
        RECT 1417.360 1576.620 1417.620 1576.880 ;
        RECT 2304.700 1576.620 2304.960 1576.880 ;
      LAYER met2 ;
        RECT 1387.360 1700.340 1387.640 1704.000 ;
        RECT 1387.360 1700.000 1387.660 1700.340 ;
        RECT 1387.520 1689.450 1387.660 1700.000 ;
        RECT 1387.460 1689.130 1387.720 1689.450 ;
        RECT 1417.360 1675.870 1417.620 1676.190 ;
        RECT 1417.420 1576.910 1417.560 1675.870 ;
        RECT 1417.360 1576.590 1417.620 1576.910 ;
        RECT 2304.700 1576.590 2304.960 1576.910 ;
        RECT 2304.760 17.410 2304.900 1576.590 ;
        RECT 2304.760 17.270 2310.420 17.410 ;
        RECT 2310.280 2.400 2310.420 17.270 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1400.845 1630.045 1401.015 1630.895 ;
        RECT 1448.685 1630.045 1448.855 1632.255 ;
        RECT 1496.985 1631.405 1497.155 1632.255 ;
        RECT 1497.445 1631.065 1497.615 1632.255 ;
        RECT 1544.825 1631.065 1544.995 1632.255 ;
        RECT 1545.745 1631.405 1545.915 1632.255 ;
        RECT 1593.585 1631.405 1593.755 1632.255 ;
        RECT 1594.045 1631.065 1594.215 1632.255 ;
        RECT 1641.885 1631.065 1642.055 1632.255 ;
        RECT 1690.645 1631.065 1690.815 1632.255 ;
        RECT 1738.025 1631.065 1738.195 1632.255 ;
        RECT 1786.785 1632.085 1786.955 1633.955 ;
      LAYER mcon ;
        RECT 1786.785 1633.785 1786.955 1633.955 ;
        RECT 1448.685 1632.085 1448.855 1632.255 ;
        RECT 1400.845 1630.725 1401.015 1630.895 ;
        RECT 1496.985 1632.085 1497.155 1632.255 ;
        RECT 1497.445 1632.085 1497.615 1632.255 ;
        RECT 1544.825 1632.085 1544.995 1632.255 ;
        RECT 1545.745 1632.085 1545.915 1632.255 ;
        RECT 1593.585 1632.085 1593.755 1632.255 ;
        RECT 1594.045 1632.085 1594.215 1632.255 ;
        RECT 1641.885 1632.085 1642.055 1632.255 ;
        RECT 1690.645 1632.085 1690.815 1632.255 ;
        RECT 1738.025 1632.085 1738.195 1632.255 ;
      LAYER met1 ;
        RECT 1389.270 1685.960 1389.590 1686.020 ;
        RECT 1396.170 1685.960 1396.490 1686.020 ;
        RECT 1389.270 1685.820 1396.490 1685.960 ;
        RECT 1389.270 1685.760 1389.590 1685.820 ;
        RECT 1396.170 1685.760 1396.490 1685.820 ;
        RECT 1738.870 1633.940 1739.190 1634.000 ;
        RECT 1786.725 1633.940 1787.015 1633.985 ;
        RECT 1738.870 1633.800 1787.015 1633.940 ;
        RECT 1738.870 1633.740 1739.190 1633.800 ;
        RECT 1786.725 1633.755 1787.015 1633.800 ;
        RECT 1448.625 1632.240 1448.915 1632.285 ;
        RECT 1496.925 1632.240 1497.215 1632.285 ;
        RECT 1497.385 1632.240 1497.675 1632.285 ;
        RECT 1448.625 1632.100 1449.300 1632.240 ;
        RECT 1448.625 1632.055 1448.915 1632.100 ;
        RECT 1449.160 1631.560 1449.300 1632.100 ;
        RECT 1496.925 1632.100 1497.675 1632.240 ;
        RECT 1496.925 1632.055 1497.215 1632.100 ;
        RECT 1497.385 1632.055 1497.675 1632.100 ;
        RECT 1544.765 1632.240 1545.055 1632.285 ;
        RECT 1545.685 1632.240 1545.975 1632.285 ;
        RECT 1544.765 1632.100 1545.975 1632.240 ;
        RECT 1544.765 1632.055 1545.055 1632.100 ;
        RECT 1545.685 1632.055 1545.975 1632.100 ;
        RECT 1593.525 1632.240 1593.815 1632.285 ;
        RECT 1593.985 1632.240 1594.275 1632.285 ;
        RECT 1593.525 1632.100 1594.275 1632.240 ;
        RECT 1593.525 1632.055 1593.815 1632.100 ;
        RECT 1593.985 1632.055 1594.275 1632.100 ;
        RECT 1641.825 1632.240 1642.115 1632.285 ;
        RECT 1690.585 1632.240 1690.875 1632.285 ;
        RECT 1641.825 1632.100 1690.875 1632.240 ;
        RECT 1641.825 1632.055 1642.115 1632.100 ;
        RECT 1690.585 1632.055 1690.875 1632.100 ;
        RECT 1737.965 1632.240 1738.255 1632.285 ;
        RECT 1738.870 1632.240 1739.190 1632.300 ;
        RECT 1737.965 1632.100 1739.190 1632.240 ;
        RECT 1737.965 1632.055 1738.255 1632.100 ;
        RECT 1738.870 1632.040 1739.190 1632.100 ;
        RECT 1786.725 1632.240 1787.015 1632.285 ;
        RECT 2325.370 1632.240 2325.690 1632.300 ;
        RECT 1786.725 1632.100 2325.690 1632.240 ;
        RECT 1786.725 1632.055 1787.015 1632.100 ;
        RECT 2325.370 1632.040 2325.690 1632.100 ;
        RECT 1496.925 1631.560 1497.215 1631.605 ;
        RECT 1449.160 1631.420 1497.215 1631.560 ;
        RECT 1496.925 1631.375 1497.215 1631.420 ;
        RECT 1545.685 1631.560 1545.975 1631.605 ;
        RECT 1593.525 1631.560 1593.815 1631.605 ;
        RECT 1545.685 1631.420 1593.815 1631.560 ;
        RECT 1545.685 1631.375 1545.975 1631.420 ;
        RECT 1593.525 1631.375 1593.815 1631.420 ;
        RECT 1497.385 1631.220 1497.675 1631.265 ;
        RECT 1544.765 1631.220 1545.055 1631.265 ;
        RECT 1497.385 1631.080 1545.055 1631.220 ;
        RECT 1497.385 1631.035 1497.675 1631.080 ;
        RECT 1544.765 1631.035 1545.055 1631.080 ;
        RECT 1593.985 1631.220 1594.275 1631.265 ;
        RECT 1641.825 1631.220 1642.115 1631.265 ;
        RECT 1593.985 1631.080 1642.115 1631.220 ;
        RECT 1593.985 1631.035 1594.275 1631.080 ;
        RECT 1641.825 1631.035 1642.115 1631.080 ;
        RECT 1690.585 1631.220 1690.875 1631.265 ;
        RECT 1737.965 1631.220 1738.255 1631.265 ;
        RECT 1690.585 1631.080 1738.255 1631.220 ;
        RECT 1690.585 1631.035 1690.875 1631.080 ;
        RECT 1737.965 1631.035 1738.255 1631.080 ;
        RECT 1396.170 1630.880 1396.490 1630.940 ;
        RECT 1400.785 1630.880 1401.075 1630.925 ;
        RECT 1396.170 1630.740 1401.075 1630.880 ;
        RECT 1396.170 1630.680 1396.490 1630.740 ;
        RECT 1400.785 1630.695 1401.075 1630.740 ;
        RECT 1400.785 1630.200 1401.075 1630.245 ;
        RECT 1448.625 1630.200 1448.915 1630.245 ;
        RECT 1400.785 1630.060 1448.915 1630.200 ;
        RECT 1400.785 1630.015 1401.075 1630.060 ;
        RECT 1448.625 1630.015 1448.915 1630.060 ;
      LAYER via ;
        RECT 1389.300 1685.760 1389.560 1686.020 ;
        RECT 1396.200 1685.760 1396.460 1686.020 ;
        RECT 1738.900 1633.740 1739.160 1634.000 ;
        RECT 1738.900 1632.040 1739.160 1632.300 ;
        RECT 2325.400 1632.040 2325.660 1632.300 ;
        RECT 1396.200 1630.680 1396.460 1630.940 ;
      LAYER met2 ;
        RECT 1389.200 1700.340 1389.480 1704.000 ;
        RECT 1389.200 1700.000 1389.500 1700.340 ;
        RECT 1389.360 1686.050 1389.500 1700.000 ;
        RECT 1389.300 1685.730 1389.560 1686.050 ;
        RECT 1396.200 1685.730 1396.460 1686.050 ;
        RECT 1396.260 1630.970 1396.400 1685.730 ;
        RECT 1738.900 1633.710 1739.160 1634.030 ;
        RECT 1738.960 1632.330 1739.100 1633.710 ;
        RECT 1738.900 1632.010 1739.160 1632.330 ;
        RECT 2325.400 1632.010 2325.660 1632.330 ;
        RECT 1396.200 1630.650 1396.460 1630.970 ;
        RECT 2325.460 17.410 2325.600 1632.010 ;
        RECT 2325.460 17.270 2328.360 17.410 ;
        RECT 2328.220 2.400 2328.360 17.270 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1391.110 1660.120 1391.430 1660.180 ;
        RECT 2339.170 1660.120 2339.490 1660.180 ;
        RECT 1391.110 1659.980 2339.490 1660.120 ;
        RECT 1391.110 1659.920 1391.430 1659.980 ;
        RECT 2339.170 1659.920 2339.490 1659.980 ;
        RECT 2339.170 17.580 2339.490 17.640 ;
        RECT 2345.610 17.580 2345.930 17.640 ;
        RECT 2339.170 17.440 2345.930 17.580 ;
        RECT 2339.170 17.380 2339.490 17.440 ;
        RECT 2345.610 17.380 2345.930 17.440 ;
      LAYER via ;
        RECT 1391.140 1659.920 1391.400 1660.180 ;
        RECT 2339.200 1659.920 2339.460 1660.180 ;
        RECT 2339.200 17.380 2339.460 17.640 ;
        RECT 2345.640 17.380 2345.900 17.640 ;
      LAYER met2 ;
        RECT 1391.040 1700.340 1391.320 1704.000 ;
        RECT 1391.040 1700.000 1391.340 1700.340 ;
        RECT 1391.200 1660.210 1391.340 1700.000 ;
        RECT 1391.140 1659.890 1391.400 1660.210 ;
        RECT 2339.200 1659.890 2339.460 1660.210 ;
        RECT 2339.260 17.670 2339.400 1659.890 ;
        RECT 2339.200 17.350 2339.460 17.670 ;
        RECT 2345.640 17.350 2345.900 17.670 ;
        RECT 2345.700 2.400 2345.840 17.350 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1386.970 1685.620 1387.290 1685.680 ;
        RECT 1392.950 1685.620 1393.270 1685.680 ;
        RECT 1386.970 1685.480 1393.270 1685.620 ;
        RECT 1386.970 1685.420 1387.290 1685.480 ;
        RECT 1392.950 1685.420 1393.270 1685.480 ;
        RECT 1386.970 1645.840 1387.290 1645.900 ;
        RECT 2359.870 1645.840 2360.190 1645.900 ;
        RECT 1386.970 1645.700 2360.190 1645.840 ;
        RECT 1386.970 1645.640 1387.290 1645.700 ;
        RECT 2359.870 1645.640 2360.190 1645.700 ;
      LAYER via ;
        RECT 1387.000 1685.420 1387.260 1685.680 ;
        RECT 1392.980 1685.420 1393.240 1685.680 ;
        RECT 1387.000 1645.640 1387.260 1645.900 ;
        RECT 2359.900 1645.640 2360.160 1645.900 ;
      LAYER met2 ;
        RECT 1392.880 1700.340 1393.160 1704.000 ;
        RECT 1392.880 1700.000 1393.180 1700.340 ;
        RECT 1393.040 1685.710 1393.180 1700.000 ;
        RECT 1387.000 1685.390 1387.260 1685.710 ;
        RECT 1392.980 1685.390 1393.240 1685.710 ;
        RECT 1387.060 1645.930 1387.200 1685.390 ;
        RECT 1387.000 1645.610 1387.260 1645.930 ;
        RECT 2359.900 1645.610 2360.160 1645.930 ;
        RECT 2359.960 16.730 2360.100 1645.610 ;
        RECT 2359.960 16.590 2363.780 16.730 ;
        RECT 2363.640 2.400 2363.780 16.590 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1394.790 1677.120 1395.110 1677.180 ;
        RECT 1397.550 1677.120 1397.870 1677.180 ;
        RECT 1394.790 1676.980 1397.870 1677.120 ;
        RECT 1394.790 1676.920 1395.110 1676.980 ;
        RECT 1397.550 1676.920 1397.870 1676.980 ;
        RECT 1396.630 1631.900 1396.950 1631.960 ;
        RECT 1397.550 1631.900 1397.870 1631.960 ;
        RECT 1396.630 1631.760 1397.870 1631.900 ;
        RECT 1396.630 1631.700 1396.950 1631.760 ;
        RECT 1397.550 1631.700 1397.870 1631.760 ;
        RECT 1396.630 1604.700 1396.950 1604.760 ;
        RECT 2380.570 1604.700 2380.890 1604.760 ;
        RECT 1396.630 1604.560 2380.890 1604.700 ;
        RECT 1396.630 1604.500 1396.950 1604.560 ;
        RECT 2380.570 1604.500 2380.890 1604.560 ;
      LAYER via ;
        RECT 1394.820 1676.920 1395.080 1677.180 ;
        RECT 1397.580 1676.920 1397.840 1677.180 ;
        RECT 1396.660 1631.700 1396.920 1631.960 ;
        RECT 1397.580 1631.700 1397.840 1631.960 ;
        RECT 1396.660 1604.500 1396.920 1604.760 ;
        RECT 2380.600 1604.500 2380.860 1604.760 ;
      LAYER met2 ;
        RECT 1394.720 1700.340 1395.000 1704.000 ;
        RECT 1394.720 1700.000 1395.020 1700.340 ;
        RECT 1394.880 1677.210 1395.020 1700.000 ;
        RECT 1394.820 1676.890 1395.080 1677.210 ;
        RECT 1397.580 1676.890 1397.840 1677.210 ;
        RECT 1397.640 1631.990 1397.780 1676.890 ;
        RECT 1396.660 1631.670 1396.920 1631.990 ;
        RECT 1397.580 1631.670 1397.840 1631.990 ;
        RECT 1396.720 1604.790 1396.860 1631.670 ;
        RECT 1396.660 1604.470 1396.920 1604.790 ;
        RECT 2380.600 1604.470 2380.860 1604.790 ;
        RECT 2380.660 16.730 2380.800 1604.470 ;
        RECT 2380.660 16.590 2381.720 16.730 ;
        RECT 2381.580 2.400 2381.720 16.590 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1397.090 1570.020 1397.410 1570.080 ;
        RECT 2394.370 1570.020 2394.690 1570.080 ;
        RECT 1397.090 1569.880 2394.690 1570.020 ;
        RECT 1397.090 1569.820 1397.410 1569.880 ;
        RECT 2394.370 1569.820 2394.690 1569.880 ;
      LAYER via ;
        RECT 1397.120 1569.820 1397.380 1570.080 ;
        RECT 2394.400 1569.820 2394.660 1570.080 ;
      LAYER met2 ;
        RECT 1396.560 1700.340 1396.840 1704.000 ;
        RECT 1396.560 1700.000 1396.860 1700.340 ;
        RECT 1396.720 1666.410 1396.860 1700.000 ;
        RECT 1396.720 1666.270 1397.320 1666.410 ;
        RECT 1397.180 1570.110 1397.320 1666.270 ;
        RECT 1397.120 1569.790 1397.380 1570.110 ;
        RECT 2394.400 1569.790 2394.660 1570.110 ;
        RECT 2394.460 16.730 2394.600 1569.790 ;
        RECT 2394.460 16.590 2399.660 16.730 ;
        RECT 2399.520 2.400 2399.660 16.590 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1214.930 1686.300 1215.250 1686.360 ;
        RECT 1231.030 1686.300 1231.350 1686.360 ;
        RECT 1214.930 1686.160 1231.350 1686.300 ;
        RECT 1214.930 1686.100 1215.250 1686.160 ;
        RECT 1231.030 1686.100 1231.350 1686.160 ;
        RECT 800.010 1673.720 800.330 1673.780 ;
        RECT 1214.930 1673.720 1215.250 1673.780 ;
        RECT 800.010 1673.580 1215.250 1673.720 ;
        RECT 800.010 1673.520 800.330 1673.580 ;
        RECT 1214.930 1673.520 1215.250 1673.580 ;
        RECT 793.570 20.980 793.890 21.040 ;
        RECT 800.010 20.980 800.330 21.040 ;
        RECT 793.570 20.840 800.330 20.980 ;
        RECT 793.570 20.780 793.890 20.840 ;
        RECT 800.010 20.780 800.330 20.840 ;
      LAYER via ;
        RECT 1214.960 1686.100 1215.220 1686.360 ;
        RECT 1231.060 1686.100 1231.320 1686.360 ;
        RECT 800.040 1673.520 800.300 1673.780 ;
        RECT 1214.960 1673.520 1215.220 1673.780 ;
        RECT 793.600 20.780 793.860 21.040 ;
        RECT 800.040 20.780 800.300 21.040 ;
      LAYER met2 ;
        RECT 1230.960 1700.340 1231.240 1704.000 ;
        RECT 1230.960 1700.000 1231.260 1700.340 ;
        RECT 1231.120 1686.390 1231.260 1700.000 ;
        RECT 1214.960 1686.070 1215.220 1686.390 ;
        RECT 1231.060 1686.070 1231.320 1686.390 ;
        RECT 1215.020 1673.810 1215.160 1686.070 ;
        RECT 800.040 1673.490 800.300 1673.810 ;
        RECT 1214.960 1673.490 1215.220 1673.810 ;
        RECT 800.100 21.070 800.240 1673.490 ;
        RECT 793.600 20.750 793.860 21.070 ;
        RECT 800.040 20.750 800.300 21.070 ;
        RECT 793.660 2.400 793.800 20.750 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 641.310 1653.320 641.630 1653.380 ;
        RECT 1215.390 1653.320 1215.710 1653.380 ;
        RECT 641.310 1653.180 1215.710 1653.320 ;
        RECT 641.310 1653.120 641.630 1653.180 ;
        RECT 1215.390 1653.120 1215.710 1653.180 ;
      LAYER via ;
        RECT 641.340 1653.120 641.600 1653.380 ;
        RECT 1215.420 1653.120 1215.680 1653.380 ;
      LAYER met2 ;
        RECT 1215.320 1700.340 1215.600 1704.000 ;
        RECT 1215.320 1700.000 1215.620 1700.340 ;
        RECT 1215.480 1653.410 1215.620 1700.000 ;
        RECT 641.340 1653.090 641.600 1653.410 ;
        RECT 1215.420 1653.090 1215.680 1653.410 ;
        RECT 641.400 17.410 641.540 1653.090 ;
        RECT 639.100 17.270 641.540 17.410 ;
        RECT 639.100 2.400 639.240 17.270 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1398.930 1632.380 1399.250 1632.640 ;
        RECT 1397.550 1631.220 1397.870 1631.280 ;
        RECT 1399.020 1631.220 1399.160 1632.380 ;
        RECT 1397.550 1631.080 1399.160 1631.220 ;
        RECT 1397.550 1631.020 1397.870 1631.080 ;
        RECT 1397.550 1563.220 1397.870 1563.280 ;
        RECT 2421.970 1563.220 2422.290 1563.280 ;
        RECT 1397.550 1563.080 2422.290 1563.220 ;
        RECT 1397.550 1563.020 1397.870 1563.080 ;
        RECT 2421.970 1563.020 2422.290 1563.080 ;
      LAYER via ;
        RECT 1398.960 1632.380 1399.220 1632.640 ;
        RECT 1397.580 1631.020 1397.840 1631.280 ;
        RECT 1397.580 1563.020 1397.840 1563.280 ;
        RECT 2422.000 1563.020 2422.260 1563.280 ;
      LAYER met2 ;
        RECT 1398.860 1700.340 1399.140 1704.000 ;
        RECT 1398.860 1700.000 1399.160 1700.340 ;
        RECT 1399.020 1632.670 1399.160 1700.000 ;
        RECT 1398.960 1632.350 1399.220 1632.670 ;
        RECT 1397.580 1630.990 1397.840 1631.310 ;
        RECT 1397.640 1563.310 1397.780 1630.990 ;
        RECT 1397.580 1562.990 1397.840 1563.310 ;
        RECT 2422.000 1562.990 2422.260 1563.310 ;
        RECT 2422.060 17.410 2422.200 1562.990 ;
        RECT 2422.060 17.270 2423.120 17.410 ;
        RECT 2422.980 2.400 2423.120 17.270 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1400.770 1683.920 1401.090 1683.980 ;
        RECT 1402.150 1683.920 1402.470 1683.980 ;
        RECT 1400.770 1683.780 1402.470 1683.920 ;
        RECT 1400.770 1683.720 1401.090 1683.780 ;
        RECT 1402.150 1683.720 1402.470 1683.780 ;
        RECT 1403.530 1597.560 1403.850 1597.620 ;
        RECT 2435.770 1597.560 2436.090 1597.620 ;
        RECT 1403.530 1597.420 2436.090 1597.560 ;
        RECT 1403.530 1597.360 1403.850 1597.420 ;
        RECT 2435.770 1597.360 2436.090 1597.420 ;
      LAYER via ;
        RECT 1400.800 1683.720 1401.060 1683.980 ;
        RECT 1402.180 1683.720 1402.440 1683.980 ;
        RECT 1403.560 1597.360 1403.820 1597.620 ;
        RECT 2435.800 1597.360 2436.060 1597.620 ;
      LAYER met2 ;
        RECT 1400.700 1700.340 1400.980 1704.000 ;
        RECT 1400.700 1700.000 1401.000 1700.340 ;
        RECT 1400.860 1684.010 1401.000 1700.000 ;
        RECT 1400.800 1683.690 1401.060 1684.010 ;
        RECT 1402.180 1683.690 1402.440 1684.010 ;
        RECT 1402.240 1677.290 1402.380 1683.690 ;
        RECT 1402.240 1677.150 1403.300 1677.290 ;
        RECT 1403.160 1631.050 1403.300 1677.150 ;
        RECT 1403.160 1630.910 1403.760 1631.050 ;
        RECT 1403.620 1597.650 1403.760 1630.910 ;
        RECT 1403.560 1597.330 1403.820 1597.650 ;
        RECT 2435.800 1597.330 2436.060 1597.650 ;
        RECT 2435.860 17.410 2436.000 1597.330 ;
        RECT 2435.860 17.270 2441.060 17.410 ;
        RECT 2440.920 2.400 2441.060 17.270 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1404.450 1556.080 1404.770 1556.140 ;
        RECT 2456.470 1556.080 2456.790 1556.140 ;
        RECT 1404.450 1555.940 2456.790 1556.080 ;
        RECT 1404.450 1555.880 1404.770 1555.940 ;
        RECT 2456.470 1555.880 2456.790 1555.940 ;
      LAYER via ;
        RECT 1404.480 1555.880 1404.740 1556.140 ;
        RECT 2456.500 1555.880 2456.760 1556.140 ;
      LAYER met2 ;
        RECT 1402.540 1700.340 1402.820 1704.000 ;
        RECT 1402.540 1700.000 1402.840 1700.340 ;
        RECT 1402.700 1677.970 1402.840 1700.000 ;
        RECT 1402.700 1677.830 1404.220 1677.970 ;
        RECT 1404.080 1632.410 1404.220 1677.830 ;
        RECT 1404.080 1632.270 1404.680 1632.410 ;
        RECT 1404.540 1556.170 1404.680 1632.270 ;
        RECT 1404.480 1555.850 1404.740 1556.170 ;
        RECT 2456.500 1555.850 2456.760 1556.170 ;
        RECT 2456.560 3.130 2456.700 1555.850 ;
        RECT 2456.560 2.990 2459.000 3.130 ;
        RECT 2458.860 2.400 2459.000 2.990 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1404.910 1549.280 1405.230 1549.340 ;
        RECT 2470.270 1549.280 2470.590 1549.340 ;
        RECT 1404.910 1549.140 2470.590 1549.280 ;
        RECT 1404.910 1549.080 1405.230 1549.140 ;
        RECT 2470.270 1549.080 2470.590 1549.140 ;
        RECT 2470.270 16.900 2470.590 16.960 ;
        RECT 2476.710 16.900 2477.030 16.960 ;
        RECT 2470.270 16.760 2477.030 16.900 ;
        RECT 2470.270 16.700 2470.590 16.760 ;
        RECT 2476.710 16.700 2477.030 16.760 ;
      LAYER via ;
        RECT 1404.940 1549.080 1405.200 1549.340 ;
        RECT 2470.300 1549.080 2470.560 1549.340 ;
        RECT 2470.300 16.700 2470.560 16.960 ;
        RECT 2476.740 16.700 2477.000 16.960 ;
      LAYER met2 ;
        RECT 1404.380 1700.340 1404.660 1704.000 ;
        RECT 1404.380 1700.000 1404.680 1700.340 ;
        RECT 1404.540 1675.250 1404.680 1700.000 ;
        RECT 1404.540 1675.110 1405.140 1675.250 ;
        RECT 1405.000 1549.370 1405.140 1675.110 ;
        RECT 1404.940 1549.050 1405.200 1549.370 ;
        RECT 2470.300 1549.050 2470.560 1549.370 ;
        RECT 2470.360 16.990 2470.500 1549.050 ;
        RECT 2470.300 16.670 2470.560 16.990 ;
        RECT 2476.740 16.670 2477.000 16.990 ;
        RECT 2476.800 2.400 2476.940 16.670 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1405.370 1542.480 1405.690 1542.540 ;
        RECT 2490.970 1542.480 2491.290 1542.540 ;
        RECT 1405.370 1542.340 2491.290 1542.480 ;
        RECT 1405.370 1542.280 1405.690 1542.340 ;
        RECT 2490.970 1542.280 2491.290 1542.340 ;
        RECT 2490.970 2.960 2491.290 3.020 ;
        RECT 2494.650 2.960 2494.970 3.020 ;
        RECT 2490.970 2.820 2494.970 2.960 ;
        RECT 2490.970 2.760 2491.290 2.820 ;
        RECT 2494.650 2.760 2494.970 2.820 ;
      LAYER via ;
        RECT 1405.400 1542.280 1405.660 1542.540 ;
        RECT 2491.000 1542.280 2491.260 1542.540 ;
        RECT 2491.000 2.760 2491.260 3.020 ;
        RECT 2494.680 2.760 2494.940 3.020 ;
      LAYER met2 ;
        RECT 1406.220 1700.340 1406.500 1704.000 ;
        RECT 1406.220 1700.000 1406.520 1700.340 ;
        RECT 1406.380 1660.970 1406.520 1700.000 ;
        RECT 1405.460 1660.830 1406.520 1660.970 ;
        RECT 1405.460 1542.570 1405.600 1660.830 ;
        RECT 1405.400 1542.250 1405.660 1542.570 ;
        RECT 2491.000 1542.250 2491.260 1542.570 ;
        RECT 2491.060 3.050 2491.200 1542.250 ;
        RECT 2491.000 2.730 2491.260 3.050 ;
        RECT 2494.680 2.730 2494.940 3.050 ;
        RECT 2494.740 2.400 2494.880 2.730 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1409.050 1625.100 1409.370 1625.160 ;
        RECT 2511.670 1625.100 2511.990 1625.160 ;
        RECT 1409.050 1624.960 2511.990 1625.100 ;
        RECT 1409.050 1624.900 1409.370 1624.960 ;
        RECT 2511.670 1624.900 2511.990 1624.960 ;
      LAYER via ;
        RECT 1409.080 1624.900 1409.340 1625.160 ;
        RECT 2511.700 1624.900 2511.960 1625.160 ;
      LAYER met2 ;
        RECT 1408.060 1700.340 1408.340 1704.000 ;
        RECT 1408.060 1700.000 1408.360 1700.340 ;
        RECT 1408.220 1656.210 1408.360 1700.000 ;
        RECT 1408.220 1656.070 1409.280 1656.210 ;
        RECT 1409.140 1625.190 1409.280 1656.070 ;
        RECT 1409.080 1624.870 1409.340 1625.190 ;
        RECT 2511.700 1624.870 2511.960 1625.190 ;
        RECT 2511.760 17.410 2511.900 1624.870 ;
        RECT 2511.760 17.270 2512.360 17.410 ;
        RECT 2512.220 2.400 2512.360 17.270 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1410.430 1631.900 1410.750 1631.960 ;
        RECT 1411.810 1631.900 1412.130 1631.960 ;
        RECT 1410.430 1631.760 1412.130 1631.900 ;
        RECT 1410.430 1631.700 1410.750 1631.760 ;
        RECT 1411.810 1631.700 1412.130 1631.760 ;
        RECT 1411.810 1590.420 1412.130 1590.480 ;
        RECT 2525.470 1590.420 2525.790 1590.480 ;
        RECT 1411.810 1590.280 2525.790 1590.420 ;
        RECT 1411.810 1590.220 1412.130 1590.280 ;
        RECT 2525.470 1590.220 2525.790 1590.280 ;
      LAYER via ;
        RECT 1410.460 1631.700 1410.720 1631.960 ;
        RECT 1411.840 1631.700 1412.100 1631.960 ;
        RECT 1411.840 1590.220 1412.100 1590.480 ;
        RECT 2525.500 1590.220 2525.760 1590.480 ;
      LAYER met2 ;
        RECT 1409.900 1700.340 1410.180 1704.000 ;
        RECT 1409.900 1700.000 1410.200 1700.340 ;
        RECT 1410.060 1668.450 1410.200 1700.000 ;
        RECT 1410.060 1668.310 1410.660 1668.450 ;
        RECT 1410.520 1631.990 1410.660 1668.310 ;
        RECT 1410.460 1631.670 1410.720 1631.990 ;
        RECT 1411.840 1631.670 1412.100 1631.990 ;
        RECT 1411.900 1590.510 1412.040 1631.670 ;
        RECT 1411.840 1590.190 1412.100 1590.510 ;
        RECT 2525.500 1590.190 2525.760 1590.510 ;
        RECT 2525.560 17.410 2525.700 1590.190 ;
        RECT 2525.560 17.270 2530.300 17.410 ;
        RECT 2530.160 2.400 2530.300 17.270 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1409.050 1685.280 1409.370 1685.340 ;
        RECT 1411.810 1685.280 1412.130 1685.340 ;
        RECT 1409.050 1685.140 1412.130 1685.280 ;
        RECT 1409.050 1685.080 1409.370 1685.140 ;
        RECT 1411.810 1685.080 1412.130 1685.140 ;
        RECT 1409.510 1639.040 1409.830 1639.100 ;
        RECT 2546.170 1639.040 2546.490 1639.100 ;
        RECT 1409.510 1638.900 2546.490 1639.040 ;
        RECT 1409.510 1638.840 1409.830 1638.900 ;
        RECT 2546.170 1638.840 2546.490 1638.900 ;
      LAYER via ;
        RECT 1409.080 1685.080 1409.340 1685.340 ;
        RECT 1411.840 1685.080 1412.100 1685.340 ;
        RECT 1409.540 1638.840 1409.800 1639.100 ;
        RECT 2546.200 1638.840 2546.460 1639.100 ;
      LAYER met2 ;
        RECT 1411.740 1700.340 1412.020 1704.000 ;
        RECT 1411.740 1700.000 1412.040 1700.340 ;
        RECT 1411.900 1685.370 1412.040 1700.000 ;
        RECT 1409.080 1685.050 1409.340 1685.370 ;
        RECT 1411.840 1685.050 1412.100 1685.370 ;
        RECT 1409.140 1667.090 1409.280 1685.050 ;
        RECT 1409.140 1666.950 1409.740 1667.090 ;
        RECT 1409.600 1639.130 1409.740 1666.950 ;
        RECT 1409.540 1638.810 1409.800 1639.130 ;
        RECT 2546.200 1638.810 2546.460 1639.130 ;
        RECT 2546.260 17.410 2546.400 1638.810 ;
        RECT 2546.260 17.270 2548.240 17.410 ;
        RECT 2548.100 2.400 2548.240 17.270 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1410.890 1683.920 1411.210 1683.980 ;
        RECT 1413.650 1683.920 1413.970 1683.980 ;
        RECT 1410.890 1683.780 1413.970 1683.920 ;
        RECT 1410.890 1683.720 1411.210 1683.780 ;
        RECT 1413.650 1683.720 1413.970 1683.780 ;
        RECT 1410.890 1535.340 1411.210 1535.400 ;
        RECT 2559.970 1535.340 2560.290 1535.400 ;
        RECT 1410.890 1535.200 2560.290 1535.340 ;
        RECT 1410.890 1535.140 1411.210 1535.200 ;
        RECT 2559.970 1535.140 2560.290 1535.200 ;
        RECT 2559.970 16.900 2560.290 16.960 ;
        RECT 2565.950 16.900 2566.270 16.960 ;
        RECT 2559.970 16.760 2566.270 16.900 ;
        RECT 2559.970 16.700 2560.290 16.760 ;
        RECT 2565.950 16.700 2566.270 16.760 ;
      LAYER via ;
        RECT 1410.920 1683.720 1411.180 1683.980 ;
        RECT 1413.680 1683.720 1413.940 1683.980 ;
        RECT 1410.920 1535.140 1411.180 1535.400 ;
        RECT 2560.000 1535.140 2560.260 1535.400 ;
        RECT 2560.000 16.700 2560.260 16.960 ;
        RECT 2565.980 16.700 2566.240 16.960 ;
      LAYER met2 ;
        RECT 1413.580 1700.340 1413.860 1704.000 ;
        RECT 1413.580 1700.000 1413.880 1700.340 ;
        RECT 1413.740 1684.010 1413.880 1700.000 ;
        RECT 1410.920 1683.690 1411.180 1684.010 ;
        RECT 1413.680 1683.690 1413.940 1684.010 ;
        RECT 1410.980 1535.430 1411.120 1683.690 ;
        RECT 1410.920 1535.110 1411.180 1535.430 ;
        RECT 2560.000 1535.110 2560.260 1535.430 ;
        RECT 2560.060 16.990 2560.200 1535.110 ;
        RECT 2560.000 16.670 2560.260 16.990 ;
        RECT 2565.980 16.670 2566.240 16.990 ;
        RECT 2566.040 2.400 2566.180 16.670 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1415.490 1683.920 1415.810 1683.980 ;
        RECT 1418.250 1683.920 1418.570 1683.980 ;
        RECT 1415.490 1683.780 1418.570 1683.920 ;
        RECT 1415.490 1683.720 1415.810 1683.780 ;
        RECT 1418.250 1683.720 1418.570 1683.780 ;
        RECT 1418.250 1583.620 1418.570 1583.680 ;
        RECT 2580.670 1583.620 2580.990 1583.680 ;
        RECT 1418.250 1583.480 2580.990 1583.620 ;
        RECT 1418.250 1583.420 1418.570 1583.480 ;
        RECT 2580.670 1583.420 2580.990 1583.480 ;
      LAYER via ;
        RECT 1415.520 1683.720 1415.780 1683.980 ;
        RECT 1418.280 1683.720 1418.540 1683.980 ;
        RECT 1418.280 1583.420 1418.540 1583.680 ;
        RECT 2580.700 1583.420 2580.960 1583.680 ;
      LAYER met2 ;
        RECT 1415.420 1700.340 1415.700 1704.000 ;
        RECT 1415.420 1700.000 1415.720 1700.340 ;
        RECT 1415.580 1684.010 1415.720 1700.000 ;
        RECT 1415.520 1683.690 1415.780 1684.010 ;
        RECT 1418.280 1683.690 1418.540 1684.010 ;
        RECT 1418.340 1583.710 1418.480 1683.690 ;
        RECT 1418.280 1583.390 1418.540 1583.710 ;
        RECT 2580.700 1583.390 2580.960 1583.710 ;
        RECT 2580.760 17.410 2580.900 1583.390 ;
        RECT 2580.760 17.270 2584.120 17.410 ;
        RECT 2583.980 2.400 2584.120 17.270 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1141.790 1685.620 1142.110 1685.680 ;
        RECT 1141.790 1685.480 1197.220 1685.620 ;
        RECT 1141.790 1685.420 1142.110 1685.480 ;
        RECT 1197.080 1685.280 1197.220 1685.480 ;
        RECT 1233.790 1685.280 1234.110 1685.340 ;
        RECT 1197.080 1685.140 1234.110 1685.280 ;
        RECT 1233.790 1685.080 1234.110 1685.140 ;
        RECT 820.710 72.320 821.030 72.380 ;
        RECT 1141.790 72.320 1142.110 72.380 ;
        RECT 820.710 72.180 1142.110 72.320 ;
        RECT 820.710 72.120 821.030 72.180 ;
        RECT 1141.790 72.120 1142.110 72.180 ;
      LAYER via ;
        RECT 1141.820 1685.420 1142.080 1685.680 ;
        RECT 1233.820 1685.080 1234.080 1685.340 ;
        RECT 820.740 72.120 821.000 72.380 ;
        RECT 1141.820 72.120 1142.080 72.380 ;
      LAYER met2 ;
        RECT 1233.720 1700.340 1234.000 1704.000 ;
        RECT 1233.720 1700.000 1234.020 1700.340 ;
        RECT 1141.820 1685.390 1142.080 1685.710 ;
        RECT 1141.880 72.410 1142.020 1685.390 ;
        RECT 1233.880 1685.370 1234.020 1700.000 ;
        RECT 1233.820 1685.050 1234.080 1685.370 ;
        RECT 820.740 72.090 821.000 72.410 ;
        RECT 1141.820 72.090 1142.080 72.410 ;
        RECT 820.800 17.410 820.940 72.090 ;
        RECT 817.580 17.270 820.940 17.410 ;
        RECT 817.580 2.400 817.720 17.270 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1417.330 1677.460 1417.650 1677.520 ;
        RECT 1420.090 1677.460 1420.410 1677.520 ;
        RECT 1417.330 1677.320 1420.410 1677.460 ;
        RECT 1417.330 1677.260 1417.650 1677.320 ;
        RECT 1420.090 1677.260 1420.410 1677.320 ;
        RECT 1420.090 1528.200 1420.410 1528.260 ;
        RECT 2601.370 1528.200 2601.690 1528.260 ;
        RECT 1420.090 1528.060 2601.690 1528.200 ;
        RECT 1420.090 1528.000 1420.410 1528.060 ;
        RECT 2601.370 1528.000 2601.690 1528.060 ;
      LAYER via ;
        RECT 1417.360 1677.260 1417.620 1677.520 ;
        RECT 1420.120 1677.260 1420.380 1677.520 ;
        RECT 1420.120 1528.000 1420.380 1528.260 ;
        RECT 2601.400 1528.000 2601.660 1528.260 ;
      LAYER met2 ;
        RECT 1417.260 1700.340 1417.540 1704.000 ;
        RECT 1417.260 1700.000 1417.560 1700.340 ;
        RECT 1417.420 1677.550 1417.560 1700.000 ;
        RECT 1417.360 1677.230 1417.620 1677.550 ;
        RECT 1420.120 1677.230 1420.380 1677.550 ;
        RECT 1420.180 1528.290 1420.320 1677.230 ;
        RECT 1420.120 1527.970 1420.380 1528.290 ;
        RECT 2601.400 1527.970 2601.660 1528.290 ;
        RECT 2601.460 2.400 2601.600 1527.970 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.170 1521.400 1419.490 1521.460 ;
        RECT 2615.170 1521.400 2615.490 1521.460 ;
        RECT 1419.170 1521.260 2615.490 1521.400 ;
        RECT 1419.170 1521.200 1419.490 1521.260 ;
        RECT 2615.170 1521.200 2615.490 1521.260 ;
      LAYER via ;
        RECT 1419.200 1521.200 1419.460 1521.460 ;
        RECT 2615.200 1521.200 2615.460 1521.460 ;
      LAYER met2 ;
        RECT 1419.100 1700.340 1419.380 1704.000 ;
        RECT 1419.100 1700.000 1419.400 1700.340 ;
        RECT 1419.260 1521.490 1419.400 1700.000 ;
        RECT 1419.200 1521.170 1419.460 1521.490 ;
        RECT 2615.200 1521.170 2615.460 1521.490 ;
        RECT 2615.260 17.410 2615.400 1521.170 ;
        RECT 2615.260 17.270 2619.540 17.410 ;
        RECT 2619.400 2.400 2619.540 17.270 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.630 1514.600 1419.950 1514.660 ;
        RECT 2635.870 1514.600 2636.190 1514.660 ;
        RECT 1419.630 1514.460 2636.190 1514.600 ;
        RECT 1419.630 1514.400 1419.950 1514.460 ;
        RECT 2635.870 1514.400 2636.190 1514.460 ;
      LAYER via ;
        RECT 1419.660 1514.400 1419.920 1514.660 ;
        RECT 2635.900 1514.400 2636.160 1514.660 ;
      LAYER met2 ;
        RECT 1420.940 1700.340 1421.220 1704.000 ;
        RECT 1420.940 1700.000 1421.240 1700.340 ;
        RECT 1421.100 1677.970 1421.240 1700.000 ;
        RECT 1419.720 1677.830 1421.240 1677.970 ;
        RECT 1419.720 1514.690 1419.860 1677.830 ;
        RECT 1419.660 1514.370 1419.920 1514.690 ;
        RECT 2635.900 1514.370 2636.160 1514.690 ;
        RECT 2635.960 17.410 2636.100 1514.370 ;
        RECT 2635.960 17.270 2637.480 17.410 ;
        RECT 2637.340 2.400 2637.480 17.270 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1422.850 1684.260 1423.170 1684.320 ;
        RECT 1425.610 1684.260 1425.930 1684.320 ;
        RECT 1422.850 1684.120 1425.930 1684.260 ;
        RECT 1422.850 1684.060 1423.170 1684.120 ;
        RECT 1425.610 1684.060 1425.930 1684.120 ;
        RECT 1425.610 1507.460 1425.930 1507.520 ;
        RECT 2649.670 1507.460 2649.990 1507.520 ;
        RECT 1425.610 1507.320 2649.990 1507.460 ;
        RECT 1425.610 1507.260 1425.930 1507.320 ;
        RECT 2649.670 1507.260 2649.990 1507.320 ;
      LAYER via ;
        RECT 1422.880 1684.060 1423.140 1684.320 ;
        RECT 1425.640 1684.060 1425.900 1684.320 ;
        RECT 1425.640 1507.260 1425.900 1507.520 ;
        RECT 2649.700 1507.260 2649.960 1507.520 ;
      LAYER met2 ;
        RECT 1422.780 1700.340 1423.060 1704.000 ;
        RECT 1422.780 1700.000 1423.080 1700.340 ;
        RECT 1422.940 1684.350 1423.080 1700.000 ;
        RECT 1422.880 1684.030 1423.140 1684.350 ;
        RECT 1425.640 1684.030 1425.900 1684.350 ;
        RECT 1425.700 1507.550 1425.840 1684.030 ;
        RECT 1425.640 1507.230 1425.900 1507.550 ;
        RECT 2649.700 1507.230 2649.960 1507.550 ;
        RECT 2649.760 17.410 2649.900 1507.230 ;
        RECT 2649.760 17.270 2655.420 17.410 ;
        RECT 2655.280 2.400 2655.420 17.270 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1424.690 1683.920 1425.010 1683.980 ;
        RECT 1426.070 1683.920 1426.390 1683.980 ;
        RECT 1424.690 1683.780 1426.390 1683.920 ;
        RECT 1424.690 1683.720 1425.010 1683.780 ;
        RECT 1426.070 1683.720 1426.390 1683.780 ;
        RECT 1426.070 1576.480 1426.390 1576.540 ;
        RECT 2670.370 1576.480 2670.690 1576.540 ;
        RECT 1426.070 1576.340 2670.690 1576.480 ;
        RECT 1426.070 1576.280 1426.390 1576.340 ;
        RECT 2670.370 1576.280 2670.690 1576.340 ;
      LAYER via ;
        RECT 1424.720 1683.720 1424.980 1683.980 ;
        RECT 1426.100 1683.720 1426.360 1683.980 ;
        RECT 1426.100 1576.280 1426.360 1576.540 ;
        RECT 2670.400 1576.280 2670.660 1576.540 ;
      LAYER met2 ;
        RECT 1424.620 1700.340 1424.900 1704.000 ;
        RECT 1424.620 1700.000 1424.920 1700.340 ;
        RECT 1424.780 1684.010 1424.920 1700.000 ;
        RECT 1424.720 1683.690 1424.980 1684.010 ;
        RECT 1426.100 1683.690 1426.360 1684.010 ;
        RECT 1426.160 1576.570 1426.300 1683.690 ;
        RECT 1426.100 1576.250 1426.360 1576.570 ;
        RECT 2670.400 1576.250 2670.660 1576.570 ;
        RECT 2670.460 17.410 2670.600 1576.250 ;
        RECT 2670.460 17.270 2672.900 17.410 ;
        RECT 2672.760 2.400 2672.900 17.270 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1422.390 1685.280 1422.710 1685.340 ;
        RECT 1426.530 1685.280 1426.850 1685.340 ;
        RECT 1422.390 1685.140 1426.850 1685.280 ;
        RECT 1422.390 1685.080 1422.710 1685.140 ;
        RECT 1426.530 1685.080 1426.850 1685.140 ;
        RECT 1422.390 1500.660 1422.710 1500.720 ;
        RECT 2684.630 1500.660 2684.950 1500.720 ;
        RECT 1422.390 1500.520 2684.950 1500.660 ;
        RECT 1422.390 1500.460 1422.710 1500.520 ;
        RECT 2684.630 1500.460 2684.950 1500.520 ;
        RECT 2684.630 18.260 2684.950 18.320 ;
        RECT 2690.610 18.260 2690.930 18.320 ;
        RECT 2684.630 18.120 2690.930 18.260 ;
        RECT 2684.630 18.060 2684.950 18.120 ;
        RECT 2690.610 18.060 2690.930 18.120 ;
      LAYER via ;
        RECT 1422.420 1685.080 1422.680 1685.340 ;
        RECT 1426.560 1685.080 1426.820 1685.340 ;
        RECT 1422.420 1500.460 1422.680 1500.720 ;
        RECT 2684.660 1500.460 2684.920 1500.720 ;
        RECT 2684.660 18.060 2684.920 18.320 ;
        RECT 2690.640 18.060 2690.900 18.320 ;
      LAYER met2 ;
        RECT 1426.460 1700.340 1426.740 1704.000 ;
        RECT 1426.460 1700.000 1426.760 1700.340 ;
        RECT 1426.620 1685.370 1426.760 1700.000 ;
        RECT 1422.420 1685.050 1422.680 1685.370 ;
        RECT 1426.560 1685.050 1426.820 1685.370 ;
        RECT 1422.480 1500.750 1422.620 1685.050 ;
        RECT 1422.420 1500.430 1422.680 1500.750 ;
        RECT 2684.660 1500.430 2684.920 1500.750 ;
        RECT 2684.720 18.350 2684.860 1500.430 ;
        RECT 2684.660 18.030 2684.920 18.350 ;
        RECT 2690.640 18.030 2690.900 18.350 ;
        RECT 2690.700 2.400 2690.840 18.030 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1428.370 1618.300 1428.690 1618.360 ;
        RECT 2704.870 1618.300 2705.190 1618.360 ;
        RECT 1428.370 1618.160 2705.190 1618.300 ;
        RECT 1428.370 1618.100 1428.690 1618.160 ;
        RECT 2704.870 1618.100 2705.190 1618.160 ;
      LAYER via ;
        RECT 1428.400 1618.100 1428.660 1618.360 ;
        RECT 2704.900 1618.100 2705.160 1618.360 ;
      LAYER met2 ;
        RECT 1428.300 1700.340 1428.580 1704.000 ;
        RECT 1428.300 1700.000 1428.600 1700.340 ;
        RECT 1428.460 1618.390 1428.600 1700.000 ;
        RECT 1428.400 1618.070 1428.660 1618.390 ;
        RECT 2704.900 1618.070 2705.160 1618.390 ;
        RECT 2704.960 17.410 2705.100 1618.070 ;
        RECT 2704.960 17.270 2708.780 17.410 ;
        RECT 2708.640 2.400 2708.780 17.270 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1430.210 1678.480 1430.530 1678.540 ;
        RECT 1431.590 1678.480 1431.910 1678.540 ;
        RECT 1430.210 1678.340 1431.910 1678.480 ;
        RECT 1430.210 1678.280 1430.530 1678.340 ;
        RECT 1431.590 1678.280 1431.910 1678.340 ;
        RECT 1432.050 1569.680 1432.370 1569.740 ;
        RECT 2725.570 1569.680 2725.890 1569.740 ;
        RECT 1432.050 1569.540 2725.890 1569.680 ;
        RECT 1432.050 1569.480 1432.370 1569.540 ;
        RECT 2725.570 1569.480 2725.890 1569.540 ;
      LAYER via ;
        RECT 1430.240 1678.280 1430.500 1678.540 ;
        RECT 1431.620 1678.280 1431.880 1678.540 ;
        RECT 1432.080 1569.480 1432.340 1569.740 ;
        RECT 2725.600 1569.480 2725.860 1569.740 ;
      LAYER met2 ;
        RECT 1430.140 1700.340 1430.420 1704.000 ;
        RECT 1430.140 1700.000 1430.440 1700.340 ;
        RECT 1430.300 1678.570 1430.440 1700.000 ;
        RECT 1430.240 1678.250 1430.500 1678.570 ;
        RECT 1431.620 1678.250 1431.880 1678.570 ;
        RECT 1431.680 1664.370 1431.820 1678.250 ;
        RECT 1431.680 1664.230 1432.280 1664.370 ;
        RECT 1432.140 1569.770 1432.280 1664.230 ;
        RECT 1432.080 1569.450 1432.340 1569.770 ;
        RECT 2725.600 1569.450 2725.860 1569.770 ;
        RECT 2725.660 17.410 2725.800 1569.450 ;
        RECT 2725.660 17.270 2726.720 17.410 ;
        RECT 2726.580 2.400 2726.720 17.270 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1432.970 1487.400 1433.290 1487.460 ;
        RECT 2739.370 1487.400 2739.690 1487.460 ;
        RECT 1432.970 1487.260 2739.690 1487.400 ;
        RECT 1432.970 1487.200 1433.290 1487.260 ;
        RECT 2739.370 1487.200 2739.690 1487.260 ;
      LAYER via ;
        RECT 1433.000 1487.200 1433.260 1487.460 ;
        RECT 2739.400 1487.200 2739.660 1487.460 ;
      LAYER met2 ;
        RECT 1431.980 1700.340 1432.260 1704.000 ;
        RECT 1431.980 1700.000 1432.280 1700.340 ;
        RECT 1432.140 1665.050 1432.280 1700.000 ;
        RECT 1432.140 1664.910 1433.200 1665.050 ;
        RECT 1433.060 1487.490 1433.200 1664.910 ;
        RECT 1433.000 1487.170 1433.260 1487.490 ;
        RECT 2739.400 1487.170 2739.660 1487.490 ;
        RECT 2739.460 17.410 2739.600 1487.170 ;
        RECT 2739.460 17.270 2744.660 17.410 ;
        RECT 2744.520 2.400 2744.660 17.270 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1433.890 1562.880 1434.210 1562.940 ;
        RECT 2760.070 1562.880 2760.390 1562.940 ;
        RECT 1433.890 1562.740 2760.390 1562.880 ;
        RECT 1433.890 1562.680 1434.210 1562.740 ;
        RECT 2760.070 1562.680 2760.390 1562.740 ;
      LAYER via ;
        RECT 1433.920 1562.680 1434.180 1562.940 ;
        RECT 2760.100 1562.680 2760.360 1562.940 ;
      LAYER met2 ;
        RECT 1433.820 1700.340 1434.100 1704.000 ;
        RECT 1433.820 1700.000 1434.120 1700.340 ;
        RECT 1433.980 1562.970 1434.120 1700.000 ;
        RECT 1433.920 1562.650 1434.180 1562.970 ;
        RECT 2760.100 1562.650 2760.360 1562.970 ;
        RECT 2760.160 17.410 2760.300 1562.650 ;
        RECT 2760.160 17.270 2762.140 17.410 ;
        RECT 2762.000 2.400 2762.140 17.270 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 841.410 1639.720 841.730 1639.780 ;
        RECT 1235.630 1639.720 1235.950 1639.780 ;
        RECT 841.410 1639.580 1235.950 1639.720 ;
        RECT 841.410 1639.520 841.730 1639.580 ;
        RECT 1235.630 1639.520 1235.950 1639.580 ;
        RECT 835.430 20.980 835.750 21.040 ;
        RECT 841.410 20.980 841.730 21.040 ;
        RECT 835.430 20.840 841.730 20.980 ;
        RECT 835.430 20.780 835.750 20.840 ;
        RECT 841.410 20.780 841.730 20.840 ;
      LAYER via ;
        RECT 841.440 1639.520 841.700 1639.780 ;
        RECT 1235.660 1639.520 1235.920 1639.780 ;
        RECT 835.460 20.780 835.720 21.040 ;
        RECT 841.440 20.780 841.700 21.040 ;
      LAYER met2 ;
        RECT 1235.560 1700.340 1235.840 1704.000 ;
        RECT 1235.560 1700.000 1235.860 1700.340 ;
        RECT 1235.720 1639.810 1235.860 1700.000 ;
        RECT 841.440 1639.490 841.700 1639.810 ;
        RECT 1235.660 1639.490 1235.920 1639.810 ;
        RECT 841.500 21.070 841.640 1639.490 ;
        RECT 835.460 20.750 835.720 21.070 ;
        RECT 841.440 20.750 841.700 21.070 ;
        RECT 835.520 2.400 835.660 20.750 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1435.730 1655.700 1436.050 1655.760 ;
        RECT 1438.490 1655.700 1438.810 1655.760 ;
        RECT 1435.730 1655.560 1438.810 1655.700 ;
        RECT 1435.730 1655.500 1436.050 1655.560 ;
        RECT 1438.490 1655.500 1438.810 1655.560 ;
        RECT 1438.490 1597.220 1438.810 1597.280 ;
        RECT 2774.330 1597.220 2774.650 1597.280 ;
        RECT 1438.490 1597.080 2774.650 1597.220 ;
        RECT 1438.490 1597.020 1438.810 1597.080 ;
        RECT 2774.330 1597.020 2774.650 1597.080 ;
      LAYER via ;
        RECT 1435.760 1655.500 1436.020 1655.760 ;
        RECT 1438.520 1655.500 1438.780 1655.760 ;
        RECT 1438.520 1597.020 1438.780 1597.280 ;
        RECT 2774.360 1597.020 2774.620 1597.280 ;
      LAYER met2 ;
        RECT 1435.660 1700.340 1435.940 1704.000 ;
        RECT 1435.660 1700.000 1435.960 1700.340 ;
        RECT 1435.820 1655.790 1435.960 1700.000 ;
        RECT 1435.760 1655.470 1436.020 1655.790 ;
        RECT 1438.520 1655.470 1438.780 1655.790 ;
        RECT 1438.580 1597.310 1438.720 1655.470 ;
        RECT 1438.520 1596.990 1438.780 1597.310 ;
        RECT 2774.360 1596.990 2774.620 1597.310 ;
        RECT 2774.420 17.410 2774.560 1596.990 ;
        RECT 2774.420 17.270 2780.080 17.410 ;
        RECT 2779.940 2.400 2780.080 17.270 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1437.110 1631.900 1437.430 1631.960 ;
        RECT 1438.950 1631.900 1439.270 1631.960 ;
        RECT 1437.110 1631.760 1439.270 1631.900 ;
        RECT 1437.110 1631.700 1437.430 1631.760 ;
        RECT 1438.950 1631.700 1439.270 1631.760 ;
        RECT 1437.110 1548.940 1437.430 1549.000 ;
        RECT 2783.990 1548.940 2784.310 1549.000 ;
        RECT 1437.110 1548.800 2784.310 1548.940 ;
        RECT 1437.110 1548.740 1437.430 1548.800 ;
        RECT 2783.990 1548.740 2784.310 1548.800 ;
        RECT 2783.990 20.640 2784.310 20.700 ;
        RECT 2797.790 20.640 2798.110 20.700 ;
        RECT 2783.990 20.500 2798.110 20.640 ;
        RECT 2783.990 20.440 2784.310 20.500 ;
        RECT 2797.790 20.440 2798.110 20.500 ;
      LAYER via ;
        RECT 1437.140 1631.700 1437.400 1631.960 ;
        RECT 1438.980 1631.700 1439.240 1631.960 ;
        RECT 1437.140 1548.740 1437.400 1549.000 ;
        RECT 2784.020 1548.740 2784.280 1549.000 ;
        RECT 2784.020 20.440 2784.280 20.700 ;
        RECT 2797.820 20.440 2798.080 20.700 ;
      LAYER met2 ;
        RECT 1437.500 1700.340 1437.780 1704.000 ;
        RECT 1437.500 1700.000 1437.800 1700.340 ;
        RECT 1437.660 1663.690 1437.800 1700.000 ;
        RECT 1437.660 1663.550 1439.180 1663.690 ;
        RECT 1439.040 1631.990 1439.180 1663.550 ;
        RECT 1437.140 1631.670 1437.400 1631.990 ;
        RECT 1438.980 1631.670 1439.240 1631.990 ;
        RECT 1437.200 1549.030 1437.340 1631.670 ;
        RECT 1437.140 1548.710 1437.400 1549.030 ;
        RECT 2784.020 1548.710 2784.280 1549.030 ;
        RECT 2784.080 20.730 2784.220 1548.710 ;
        RECT 2784.020 20.410 2784.280 20.730 ;
        RECT 2797.820 20.410 2798.080 20.730 ;
        RECT 2797.880 2.400 2798.020 20.410 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1439.410 1479.920 1439.730 1479.980 ;
        RECT 2815.270 1479.920 2815.590 1479.980 ;
        RECT 1439.410 1479.780 2815.590 1479.920 ;
        RECT 1439.410 1479.720 1439.730 1479.780 ;
        RECT 2815.270 1479.720 2815.590 1479.780 ;
      LAYER via ;
        RECT 1439.440 1479.720 1439.700 1479.980 ;
        RECT 2815.300 1479.720 2815.560 1479.980 ;
      LAYER met2 ;
        RECT 1439.340 1700.340 1439.620 1704.000 ;
        RECT 1439.340 1700.000 1439.640 1700.340 ;
        RECT 1439.500 1480.010 1439.640 1700.000 ;
        RECT 1439.440 1479.690 1439.700 1480.010 ;
        RECT 2815.300 1479.690 2815.560 1480.010 ;
        RECT 2815.360 17.410 2815.500 1479.690 ;
        RECT 2815.360 17.270 2815.960 17.410 ;
        RECT 2815.820 2.400 2815.960 17.270 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1439.870 1614.560 1440.190 1614.620 ;
        RECT 1441.250 1614.560 1441.570 1614.620 ;
        RECT 1439.870 1614.420 1441.570 1614.560 ;
        RECT 1439.870 1614.360 1440.190 1614.420 ;
        RECT 1441.250 1614.360 1441.570 1614.420 ;
        RECT 1439.870 1473.120 1440.190 1473.180 ;
        RECT 2804.690 1473.120 2805.010 1473.180 ;
        RECT 1439.870 1472.980 2805.010 1473.120 ;
        RECT 1439.870 1472.920 1440.190 1472.980 ;
        RECT 2804.690 1472.920 2805.010 1472.980 ;
        RECT 2804.690 15.200 2805.010 15.260 ;
        RECT 2833.670 15.200 2833.990 15.260 ;
        RECT 2804.690 15.060 2833.990 15.200 ;
        RECT 2804.690 15.000 2805.010 15.060 ;
        RECT 2833.670 15.000 2833.990 15.060 ;
      LAYER via ;
        RECT 1439.900 1614.360 1440.160 1614.620 ;
        RECT 1441.280 1614.360 1441.540 1614.620 ;
        RECT 1439.900 1472.920 1440.160 1473.180 ;
        RECT 2804.720 1472.920 2804.980 1473.180 ;
        RECT 2804.720 15.000 2804.980 15.260 ;
        RECT 2833.700 15.000 2833.960 15.260 ;
      LAYER met2 ;
        RECT 1441.180 1700.340 1441.460 1704.000 ;
        RECT 1441.180 1700.000 1441.480 1700.340 ;
        RECT 1441.340 1614.650 1441.480 1700.000 ;
        RECT 1439.900 1614.330 1440.160 1614.650 ;
        RECT 1441.280 1614.330 1441.540 1614.650 ;
        RECT 1439.960 1473.210 1440.100 1614.330 ;
        RECT 1439.900 1472.890 1440.160 1473.210 ;
        RECT 2804.720 1472.890 2804.980 1473.210 ;
        RECT 2804.780 15.290 2804.920 1472.890 ;
        RECT 2804.720 14.970 2804.980 15.290 ;
        RECT 2833.700 14.970 2833.960 15.290 ;
        RECT 2833.760 2.400 2833.900 14.970 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1443.090 1677.460 1443.410 1677.520 ;
        RECT 1446.310 1677.460 1446.630 1677.520 ;
        RECT 1443.090 1677.320 1446.630 1677.460 ;
        RECT 1443.090 1677.260 1443.410 1677.320 ;
        RECT 1446.310 1677.260 1446.630 1677.320 ;
        RECT 1446.310 1611.160 1446.630 1611.220 ;
        RECT 2839.190 1611.160 2839.510 1611.220 ;
        RECT 1446.310 1611.020 2839.510 1611.160 ;
        RECT 1446.310 1610.960 1446.630 1611.020 ;
        RECT 2839.190 1610.960 2839.510 1611.020 ;
        RECT 2839.190 17.920 2839.510 17.980 ;
        RECT 2851.150 17.920 2851.470 17.980 ;
        RECT 2839.190 17.780 2851.470 17.920 ;
        RECT 2839.190 17.720 2839.510 17.780 ;
        RECT 2851.150 17.720 2851.470 17.780 ;
      LAYER via ;
        RECT 1443.120 1677.260 1443.380 1677.520 ;
        RECT 1446.340 1677.260 1446.600 1677.520 ;
        RECT 1446.340 1610.960 1446.600 1611.220 ;
        RECT 2839.220 1610.960 2839.480 1611.220 ;
        RECT 2839.220 17.720 2839.480 17.980 ;
        RECT 2851.180 17.720 2851.440 17.980 ;
      LAYER met2 ;
        RECT 1443.020 1700.340 1443.300 1704.000 ;
        RECT 1443.020 1700.000 1443.320 1700.340 ;
        RECT 1443.180 1677.550 1443.320 1700.000 ;
        RECT 1443.120 1677.230 1443.380 1677.550 ;
        RECT 1446.340 1677.230 1446.600 1677.550 ;
        RECT 1446.400 1611.250 1446.540 1677.230 ;
        RECT 1446.340 1610.930 1446.600 1611.250 ;
        RECT 2839.220 1610.930 2839.480 1611.250 ;
        RECT 2839.280 18.010 2839.420 1610.930 ;
        RECT 2839.220 17.690 2839.480 18.010 ;
        RECT 2851.180 17.690 2851.440 18.010 ;
        RECT 2851.240 2.400 2851.380 17.690 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1444.930 1684.600 1445.250 1684.660 ;
        RECT 1460.110 1684.600 1460.430 1684.660 ;
        RECT 1444.930 1684.460 1460.430 1684.600 ;
        RECT 1444.930 1684.400 1445.250 1684.460 ;
        RECT 1460.110 1684.400 1460.430 1684.460 ;
        RECT 1460.110 1466.320 1460.430 1466.380 ;
        RECT 2863.570 1466.320 2863.890 1466.380 ;
        RECT 1460.110 1466.180 2863.890 1466.320 ;
        RECT 1460.110 1466.120 1460.430 1466.180 ;
        RECT 2863.570 1466.120 2863.890 1466.180 ;
      LAYER via ;
        RECT 1444.960 1684.400 1445.220 1684.660 ;
        RECT 1460.140 1684.400 1460.400 1684.660 ;
        RECT 1460.140 1466.120 1460.400 1466.380 ;
        RECT 2863.600 1466.120 2863.860 1466.380 ;
      LAYER met2 ;
        RECT 1444.860 1700.340 1445.140 1704.000 ;
        RECT 1444.860 1700.000 1445.160 1700.340 ;
        RECT 1445.020 1684.690 1445.160 1700.000 ;
        RECT 1444.960 1684.370 1445.220 1684.690 ;
        RECT 1460.140 1684.370 1460.400 1684.690 ;
        RECT 1460.200 1466.410 1460.340 1684.370 ;
        RECT 1460.140 1466.090 1460.400 1466.410 ;
        RECT 2863.600 1466.090 2863.860 1466.410 ;
        RECT 2863.660 16.730 2863.800 1466.090 ;
        RECT 2863.660 16.590 2869.320 16.730 ;
        RECT 2869.180 2.400 2869.320 16.590 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1443.165 1647.725 1443.335 1678.495 ;
      LAYER mcon ;
        RECT 1443.165 1678.325 1443.335 1678.495 ;
      LAYER met1 ;
        RECT 1443.105 1678.480 1443.395 1678.525 ;
        RECT 1446.770 1678.480 1447.090 1678.540 ;
        RECT 1443.105 1678.340 1447.090 1678.480 ;
        RECT 1443.105 1678.295 1443.395 1678.340 ;
        RECT 1446.770 1678.280 1447.090 1678.340 ;
        RECT 1443.090 1647.880 1443.410 1647.940 ;
        RECT 1442.895 1647.740 1443.410 1647.880 ;
        RECT 1443.090 1647.680 1443.410 1647.740 ;
        RECT 1443.090 1542.140 1443.410 1542.200 ;
        RECT 2874.150 1542.140 2874.470 1542.200 ;
        RECT 1443.090 1542.000 2874.470 1542.140 ;
        RECT 1443.090 1541.940 1443.410 1542.000 ;
        RECT 2874.150 1541.940 2874.470 1542.000 ;
        RECT 2874.150 16.560 2874.470 16.620 ;
        RECT 2887.030 16.560 2887.350 16.620 ;
        RECT 2874.150 16.420 2887.350 16.560 ;
        RECT 2874.150 16.360 2874.470 16.420 ;
        RECT 2887.030 16.360 2887.350 16.420 ;
      LAYER via ;
        RECT 1446.800 1678.280 1447.060 1678.540 ;
        RECT 1443.120 1647.680 1443.380 1647.940 ;
        RECT 1443.120 1541.940 1443.380 1542.200 ;
        RECT 2874.180 1541.940 2874.440 1542.200 ;
        RECT 2874.180 16.360 2874.440 16.620 ;
        RECT 2887.060 16.360 2887.320 16.620 ;
      LAYER met2 ;
        RECT 1446.700 1700.340 1446.980 1704.000 ;
        RECT 1446.700 1700.000 1447.000 1700.340 ;
        RECT 1446.860 1678.570 1447.000 1700.000 ;
        RECT 1446.800 1678.250 1447.060 1678.570 ;
        RECT 1443.120 1647.650 1443.380 1647.970 ;
        RECT 1443.180 1542.230 1443.320 1647.650 ;
        RECT 1443.120 1541.910 1443.380 1542.230 ;
        RECT 2874.180 1541.910 2874.440 1542.230 ;
        RECT 2874.240 16.650 2874.380 1541.910 ;
        RECT 2874.180 16.330 2874.440 16.650 ;
        RECT 2887.060 16.330 2887.320 16.650 ;
        RECT 2887.120 2.400 2887.260 16.330 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1447.230 1555.740 1447.550 1555.800 ;
        RECT 2859.890 1555.740 2860.210 1555.800 ;
        RECT 1447.230 1555.600 2860.210 1555.740 ;
        RECT 1447.230 1555.540 1447.550 1555.600 ;
        RECT 2859.890 1555.540 2860.210 1555.600 ;
        RECT 2859.890 18.260 2860.210 18.320 ;
        RECT 2904.970 18.260 2905.290 18.320 ;
        RECT 2859.890 18.120 2905.290 18.260 ;
        RECT 2859.890 18.060 2860.210 18.120 ;
        RECT 2904.970 18.060 2905.290 18.120 ;
      LAYER via ;
        RECT 1447.260 1555.540 1447.520 1555.800 ;
        RECT 2859.920 1555.540 2860.180 1555.800 ;
        RECT 2859.920 18.060 2860.180 18.320 ;
        RECT 2905.000 18.060 2905.260 18.320 ;
      LAYER met2 ;
        RECT 1448.540 1700.340 1448.820 1704.000 ;
        RECT 1448.540 1700.000 1448.840 1700.340 ;
        RECT 1448.700 1642.610 1448.840 1700.000 ;
        RECT 1448.240 1642.470 1448.840 1642.610 ;
        RECT 1448.240 1617.450 1448.380 1642.470 ;
        RECT 1447.320 1617.310 1448.380 1617.450 ;
        RECT 1447.320 1555.830 1447.460 1617.310 ;
        RECT 1447.260 1555.510 1447.520 1555.830 ;
        RECT 2859.920 1555.510 2860.180 1555.830 ;
        RECT 2859.980 18.350 2860.120 1555.510 ;
        RECT 2859.920 18.030 2860.180 18.350 ;
        RECT 2905.000 18.030 2905.260 18.350 ;
        RECT 2905.060 2.400 2905.200 18.030 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 855.210 1632.920 855.530 1632.980 ;
        RECT 1237.930 1632.920 1238.250 1632.980 ;
        RECT 855.210 1632.780 1238.250 1632.920 ;
        RECT 855.210 1632.720 855.530 1632.780 ;
        RECT 1237.930 1632.720 1238.250 1632.780 ;
      LAYER via ;
        RECT 855.240 1632.720 855.500 1632.980 ;
        RECT 1237.960 1632.720 1238.220 1632.980 ;
      LAYER met2 ;
        RECT 1237.400 1700.340 1237.680 1704.000 ;
        RECT 1237.400 1700.000 1237.700 1700.340 ;
        RECT 1237.560 1668.450 1237.700 1700.000 ;
        RECT 1237.560 1668.310 1238.160 1668.450 ;
        RECT 1238.020 1633.010 1238.160 1668.310 ;
        RECT 855.240 1632.690 855.500 1633.010 ;
        RECT 1237.960 1632.690 1238.220 1633.010 ;
        RECT 855.300 17.410 855.440 1632.690 ;
        RECT 853.000 17.270 855.440 17.410 ;
        RECT 853.000 2.400 853.140 17.270 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 870.850 31.860 871.170 31.920 ;
        RECT 1238.850 31.860 1239.170 31.920 ;
        RECT 870.850 31.720 1239.170 31.860 ;
        RECT 870.850 31.660 871.170 31.720 ;
        RECT 1238.850 31.660 1239.170 31.720 ;
      LAYER via ;
        RECT 870.880 31.660 871.140 31.920 ;
        RECT 1238.880 31.660 1239.140 31.920 ;
      LAYER met2 ;
        RECT 1239.240 1700.410 1239.520 1704.000 ;
        RECT 1238.940 1700.270 1239.520 1700.410 ;
        RECT 1238.940 31.950 1239.080 1700.270 ;
        RECT 1239.240 1700.000 1239.520 1700.270 ;
        RECT 870.880 31.630 871.140 31.950 ;
        RECT 1238.880 31.630 1239.140 31.950 ;
        RECT 870.940 2.400 871.080 31.630 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 888.790 32.200 889.110 32.260 ;
        RECT 1240.690 32.200 1241.010 32.260 ;
        RECT 888.790 32.060 1241.010 32.200 ;
        RECT 888.790 32.000 889.110 32.060 ;
        RECT 1240.690 32.000 1241.010 32.060 ;
      LAYER via ;
        RECT 888.820 32.000 889.080 32.260 ;
        RECT 1240.720 32.000 1240.980 32.260 ;
      LAYER met2 ;
        RECT 1241.080 1700.410 1241.360 1704.000 ;
        RECT 1240.780 1700.270 1241.360 1700.410 ;
        RECT 1240.780 32.290 1240.920 1700.270 ;
        RECT 1241.080 1700.000 1241.360 1700.270 ;
        RECT 888.820 31.970 889.080 32.290 ;
        RECT 1240.720 31.970 1240.980 32.290 ;
        RECT 888.880 2.400 889.020 31.970 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 906.730 32.540 907.050 32.600 ;
        RECT 1242.990 32.540 1243.310 32.600 ;
        RECT 906.730 32.400 1243.310 32.540 ;
        RECT 906.730 32.340 907.050 32.400 ;
        RECT 1242.990 32.340 1243.310 32.400 ;
      LAYER via ;
        RECT 906.760 32.340 907.020 32.600 ;
        RECT 1243.020 32.340 1243.280 32.600 ;
      LAYER met2 ;
        RECT 1242.920 1700.340 1243.200 1704.000 ;
        RECT 1242.920 1700.000 1243.220 1700.340 ;
        RECT 1243.080 32.630 1243.220 1700.000 ;
        RECT 906.760 32.310 907.020 32.630 ;
        RECT 1243.020 32.310 1243.280 32.630 ;
        RECT 906.820 2.400 906.960 32.310 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1244.370 1678.620 1244.690 1678.880 ;
        RECT 1244.460 1678.200 1244.600 1678.620 ;
        RECT 1244.370 1677.940 1244.690 1678.200 ;
        RECT 924.210 32.880 924.530 32.940 ;
        RECT 1244.370 32.880 1244.690 32.940 ;
        RECT 924.210 32.740 1244.690 32.880 ;
        RECT 924.210 32.680 924.530 32.740 ;
        RECT 1244.370 32.680 1244.690 32.740 ;
      LAYER via ;
        RECT 1244.400 1678.620 1244.660 1678.880 ;
        RECT 1244.400 1677.940 1244.660 1678.200 ;
        RECT 924.240 32.680 924.500 32.940 ;
        RECT 1244.400 32.680 1244.660 32.940 ;
      LAYER met2 ;
        RECT 1244.760 1700.410 1245.040 1704.000 ;
        RECT 1244.460 1700.270 1245.040 1700.410 ;
        RECT 1244.460 1678.910 1244.600 1700.270 ;
        RECT 1244.760 1700.000 1245.040 1700.270 ;
        RECT 1244.400 1678.590 1244.660 1678.910 ;
        RECT 1244.400 1677.910 1244.660 1678.230 ;
        RECT 1244.460 32.970 1244.600 1677.910 ;
        RECT 924.240 32.650 924.500 32.970 ;
        RECT 1244.400 32.650 1244.660 32.970 ;
        RECT 924.300 2.400 924.440 32.650 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 942.150 33.220 942.470 33.280 ;
        RECT 1246.670 33.220 1246.990 33.280 ;
        RECT 942.150 33.080 1246.990 33.220 ;
        RECT 942.150 33.020 942.470 33.080 ;
        RECT 1246.670 33.020 1246.990 33.080 ;
      LAYER via ;
        RECT 942.180 33.020 942.440 33.280 ;
        RECT 1246.700 33.020 1246.960 33.280 ;
      LAYER met2 ;
        RECT 1246.600 1700.340 1246.880 1704.000 ;
        RECT 1246.600 1700.000 1246.900 1700.340 ;
        RECT 1246.760 33.310 1246.900 1700.000 ;
        RECT 942.180 32.990 942.440 33.310 ;
        RECT 1246.700 32.990 1246.960 33.310 ;
        RECT 942.240 2.400 942.380 32.990 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 960.090 33.560 960.410 33.620 ;
        RECT 1248.510 33.560 1248.830 33.620 ;
        RECT 960.090 33.420 1248.830 33.560 ;
        RECT 960.090 33.360 960.410 33.420 ;
        RECT 1248.510 33.360 1248.830 33.420 ;
      LAYER via ;
        RECT 960.120 33.360 960.380 33.620 ;
        RECT 1248.540 33.360 1248.800 33.620 ;
      LAYER met2 ;
        RECT 1248.440 1700.340 1248.720 1704.000 ;
        RECT 1248.440 1700.000 1248.740 1700.340 ;
        RECT 1248.600 33.650 1248.740 1700.000 ;
        RECT 960.120 33.330 960.380 33.650 ;
        RECT 1248.540 33.330 1248.800 33.650 ;
        RECT 960.180 2.400 960.320 33.330 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 978.030 33.900 978.350 33.960 ;
        RECT 1250.350 33.900 1250.670 33.960 ;
        RECT 978.030 33.760 1250.670 33.900 ;
        RECT 978.030 33.700 978.350 33.760 ;
        RECT 1250.350 33.700 1250.670 33.760 ;
      LAYER via ;
        RECT 978.060 33.700 978.320 33.960 ;
        RECT 1250.380 33.700 1250.640 33.960 ;
      LAYER met2 ;
        RECT 1250.280 1700.340 1250.560 1704.000 ;
        RECT 1250.280 1700.000 1250.580 1700.340 ;
        RECT 1250.440 33.990 1250.580 1700.000 ;
        RECT 978.060 33.670 978.320 33.990 ;
        RECT 1250.380 33.670 1250.640 33.990 ;
        RECT 978.120 2.400 978.260 33.670 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1216.310 1678.140 1216.630 1678.200 ;
        RECT 1217.230 1678.140 1217.550 1678.200 ;
        RECT 1216.310 1678.000 1217.550 1678.140 ;
        RECT 1216.310 1677.940 1216.630 1678.000 ;
        RECT 1217.230 1677.940 1217.550 1678.000 ;
        RECT 656.950 31.180 657.270 31.240 ;
        RECT 1216.310 31.180 1216.630 31.240 ;
        RECT 656.950 31.040 1216.630 31.180 ;
        RECT 656.950 30.980 657.270 31.040 ;
        RECT 1216.310 30.980 1216.630 31.040 ;
      LAYER via ;
        RECT 1216.340 1677.940 1216.600 1678.200 ;
        RECT 1217.260 1677.940 1217.520 1678.200 ;
        RECT 656.980 30.980 657.240 31.240 ;
        RECT 1216.340 30.980 1216.600 31.240 ;
      LAYER met2 ;
        RECT 1217.160 1700.340 1217.440 1704.000 ;
        RECT 1217.160 1700.000 1217.460 1700.340 ;
        RECT 1217.320 1678.230 1217.460 1700.000 ;
        RECT 1216.340 1677.910 1216.600 1678.230 ;
        RECT 1217.260 1677.910 1217.520 1678.230 ;
        RECT 1216.400 31.270 1216.540 1677.910 ;
        RECT 656.980 30.950 657.240 31.270 ;
        RECT 1216.340 30.950 1216.600 31.270 ;
        RECT 657.040 2.400 657.180 30.950 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 995.970 34.240 996.290 34.300 ;
        RECT 1251.730 34.240 1252.050 34.300 ;
        RECT 995.970 34.100 1252.050 34.240 ;
        RECT 995.970 34.040 996.290 34.100 ;
        RECT 1251.730 34.040 1252.050 34.100 ;
      LAYER via ;
        RECT 996.000 34.040 996.260 34.300 ;
        RECT 1251.760 34.040 1252.020 34.300 ;
      LAYER met2 ;
        RECT 1252.120 1700.410 1252.400 1704.000 ;
        RECT 1251.820 1700.270 1252.400 1700.410 ;
        RECT 1251.820 34.330 1251.960 1700.270 ;
        RECT 1252.120 1700.000 1252.400 1700.270 ;
        RECT 996.000 34.010 996.260 34.330 ;
        RECT 1251.760 34.010 1252.020 34.330 ;
        RECT 996.060 2.400 996.200 34.010 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.450 30.500 1013.770 30.560 ;
        RECT 1254.030 30.500 1254.350 30.560 ;
        RECT 1013.450 30.360 1254.350 30.500 ;
        RECT 1013.450 30.300 1013.770 30.360 ;
        RECT 1254.030 30.300 1254.350 30.360 ;
      LAYER via ;
        RECT 1013.480 30.300 1013.740 30.560 ;
        RECT 1254.060 30.300 1254.320 30.560 ;
      LAYER met2 ;
        RECT 1253.960 1700.340 1254.240 1704.000 ;
        RECT 1253.960 1700.000 1254.260 1700.340 ;
        RECT 1254.120 30.590 1254.260 1700.000 ;
        RECT 1013.480 30.270 1013.740 30.590 ;
        RECT 1254.060 30.270 1254.320 30.590 ;
        RECT 1013.540 2.400 1013.680 30.270 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1255.870 1678.140 1256.190 1678.200 ;
        RECT 1257.710 1678.140 1258.030 1678.200 ;
        RECT 1255.870 1678.000 1258.030 1678.140 ;
        RECT 1255.870 1677.940 1256.190 1678.000 ;
        RECT 1257.710 1677.940 1258.030 1678.000 ;
        RECT 1034.610 1646.860 1034.930 1646.920 ;
        RECT 1257.710 1646.860 1258.030 1646.920 ;
        RECT 1034.610 1646.720 1258.030 1646.860 ;
        RECT 1034.610 1646.660 1034.930 1646.720 ;
        RECT 1257.710 1646.660 1258.030 1646.720 ;
        RECT 1031.390 2.960 1031.710 3.020 ;
        RECT 1034.610 2.960 1034.930 3.020 ;
        RECT 1031.390 2.820 1034.930 2.960 ;
        RECT 1031.390 2.760 1031.710 2.820 ;
        RECT 1034.610 2.760 1034.930 2.820 ;
      LAYER via ;
        RECT 1255.900 1677.940 1256.160 1678.200 ;
        RECT 1257.740 1677.940 1258.000 1678.200 ;
        RECT 1034.640 1646.660 1034.900 1646.920 ;
        RECT 1257.740 1646.660 1258.000 1646.920 ;
        RECT 1031.420 2.760 1031.680 3.020 ;
        RECT 1034.640 2.760 1034.900 3.020 ;
      LAYER met2 ;
        RECT 1255.800 1700.340 1256.080 1704.000 ;
        RECT 1255.800 1700.000 1256.100 1700.340 ;
        RECT 1255.960 1678.230 1256.100 1700.000 ;
        RECT 1255.900 1677.910 1256.160 1678.230 ;
        RECT 1257.740 1677.910 1258.000 1678.230 ;
        RECT 1257.800 1646.950 1257.940 1677.910 ;
        RECT 1034.640 1646.630 1034.900 1646.950 ;
        RECT 1257.740 1646.630 1258.000 1646.950 ;
        RECT 1034.700 3.050 1034.840 1646.630 ;
        RECT 1031.420 2.730 1031.680 3.050 ;
        RECT 1034.640 2.730 1034.900 3.050 ;
        RECT 1031.480 2.400 1031.620 2.730 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1055.310 1661.140 1055.630 1661.200 ;
        RECT 1256.790 1661.140 1257.110 1661.200 ;
        RECT 1055.310 1661.000 1257.110 1661.140 ;
        RECT 1055.310 1660.940 1055.630 1661.000 ;
        RECT 1256.790 1660.940 1257.110 1661.000 ;
        RECT 1049.330 20.980 1049.650 21.040 ;
        RECT 1055.310 20.980 1055.630 21.040 ;
        RECT 1049.330 20.840 1055.630 20.980 ;
        RECT 1049.330 20.780 1049.650 20.840 ;
        RECT 1055.310 20.780 1055.630 20.840 ;
      LAYER via ;
        RECT 1055.340 1660.940 1055.600 1661.200 ;
        RECT 1256.820 1660.940 1257.080 1661.200 ;
        RECT 1049.360 20.780 1049.620 21.040 ;
        RECT 1055.340 20.780 1055.600 21.040 ;
      LAYER met2 ;
        RECT 1257.640 1700.410 1257.920 1704.000 ;
        RECT 1257.340 1700.270 1257.920 1700.410 ;
        RECT 1257.340 1678.650 1257.480 1700.270 ;
        RECT 1257.640 1700.000 1257.920 1700.270 ;
        RECT 1256.880 1678.510 1257.480 1678.650 ;
        RECT 1256.880 1661.230 1257.020 1678.510 ;
        RECT 1055.340 1660.910 1055.600 1661.230 ;
        RECT 1256.820 1660.910 1257.080 1661.230 ;
        RECT 1055.400 21.070 1055.540 1660.910 ;
        RECT 1049.360 20.750 1049.620 21.070 ;
        RECT 1055.340 20.750 1055.600 21.070 ;
        RECT 1049.420 2.400 1049.560 20.750 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1257.250 1677.460 1257.570 1677.520 ;
        RECT 1258.630 1677.460 1258.950 1677.520 ;
        RECT 1257.250 1677.320 1258.950 1677.460 ;
        RECT 1257.250 1677.260 1257.570 1677.320 ;
        RECT 1258.630 1677.260 1258.950 1677.320 ;
        RECT 1069.110 1625.780 1069.430 1625.840 ;
        RECT 1257.250 1625.780 1257.570 1625.840 ;
        RECT 1069.110 1625.640 1257.570 1625.780 ;
        RECT 1069.110 1625.580 1069.430 1625.640 ;
        RECT 1257.250 1625.580 1257.570 1625.640 ;
      LAYER via ;
        RECT 1257.280 1677.260 1257.540 1677.520 ;
        RECT 1258.660 1677.260 1258.920 1677.520 ;
        RECT 1069.140 1625.580 1069.400 1625.840 ;
        RECT 1257.280 1625.580 1257.540 1625.840 ;
      LAYER met2 ;
        RECT 1259.480 1700.410 1259.760 1704.000 ;
        RECT 1259.180 1700.270 1259.760 1700.410 ;
        RECT 1259.180 1679.330 1259.320 1700.270 ;
        RECT 1259.480 1700.000 1259.760 1700.270 ;
        RECT 1258.720 1679.190 1259.320 1679.330 ;
        RECT 1258.720 1677.550 1258.860 1679.190 ;
        RECT 1257.280 1677.230 1257.540 1677.550 ;
        RECT 1258.660 1677.230 1258.920 1677.550 ;
        RECT 1257.340 1625.870 1257.480 1677.230 ;
        RECT 1069.140 1625.550 1069.400 1625.870 ;
        RECT 1257.280 1625.550 1257.540 1625.870 ;
        RECT 1069.200 18.090 1069.340 1625.550 ;
        RECT 1067.360 17.950 1069.340 18.090 ;
        RECT 1067.360 2.400 1067.500 17.950 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1089.810 1618.980 1090.130 1619.040 ;
        RECT 1261.850 1618.980 1262.170 1619.040 ;
        RECT 1089.810 1618.840 1262.170 1618.980 ;
        RECT 1089.810 1618.780 1090.130 1618.840 ;
        RECT 1261.850 1618.780 1262.170 1618.840 ;
      LAYER via ;
        RECT 1089.840 1618.780 1090.100 1619.040 ;
        RECT 1261.880 1618.780 1262.140 1619.040 ;
      LAYER met2 ;
        RECT 1261.320 1700.340 1261.600 1704.000 ;
        RECT 1261.320 1700.000 1261.620 1700.340 ;
        RECT 1261.480 1669.130 1261.620 1700.000 ;
        RECT 1261.480 1668.990 1262.080 1669.130 ;
        RECT 1261.940 1619.070 1262.080 1668.990 ;
        RECT 1089.840 1618.750 1090.100 1619.070 ;
        RECT 1261.880 1618.750 1262.140 1619.070 ;
        RECT 1089.900 18.090 1090.040 1618.750 ;
        RECT 1085.300 17.950 1090.040 18.090 ;
        RECT 1085.300 2.400 1085.440 17.950 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1263.230 1668.960 1263.550 1669.020 ;
        RECT 1236.180 1668.820 1263.550 1668.960 ;
        RECT 1103.610 1668.280 1103.930 1668.340 ;
        RECT 1236.180 1668.280 1236.320 1668.820 ;
        RECT 1263.230 1668.760 1263.550 1668.820 ;
        RECT 1103.610 1668.140 1236.320 1668.280 ;
        RECT 1103.610 1668.080 1103.930 1668.140 ;
      LAYER via ;
        RECT 1103.640 1668.080 1103.900 1668.340 ;
        RECT 1263.260 1668.760 1263.520 1669.020 ;
      LAYER met2 ;
        RECT 1263.160 1700.340 1263.440 1704.000 ;
        RECT 1263.160 1700.000 1263.460 1700.340 ;
        RECT 1263.320 1669.050 1263.460 1700.000 ;
        RECT 1263.260 1668.730 1263.520 1669.050 ;
        RECT 1103.640 1668.050 1103.900 1668.370 ;
        RECT 1103.700 16.730 1103.840 1668.050 ;
        RECT 1102.780 16.590 1103.840 16.730 ;
        RECT 1102.780 2.400 1102.920 16.590 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1234.710 1685.280 1235.030 1685.340 ;
        RECT 1264.610 1685.280 1264.930 1685.340 ;
        RECT 1234.710 1685.140 1264.930 1685.280 ;
        RECT 1234.710 1685.080 1235.030 1685.140 ;
        RECT 1264.610 1685.080 1264.930 1685.140 ;
        RECT 1124.310 1675.420 1124.630 1675.480 ;
        RECT 1234.710 1675.420 1235.030 1675.480 ;
        RECT 1124.310 1675.280 1235.030 1675.420 ;
        RECT 1124.310 1675.220 1124.630 1675.280 ;
        RECT 1234.710 1675.220 1235.030 1675.280 ;
      LAYER via ;
        RECT 1234.740 1685.080 1235.000 1685.340 ;
        RECT 1264.640 1685.080 1264.900 1685.340 ;
        RECT 1124.340 1675.220 1124.600 1675.480 ;
        RECT 1234.740 1675.220 1235.000 1675.480 ;
      LAYER met2 ;
        RECT 1265.000 1700.410 1265.280 1704.000 ;
        RECT 1264.700 1700.270 1265.280 1700.410 ;
        RECT 1264.700 1685.370 1264.840 1700.270 ;
        RECT 1265.000 1700.000 1265.280 1700.270 ;
        RECT 1234.740 1685.050 1235.000 1685.370 ;
        RECT 1264.640 1685.050 1264.900 1685.370 ;
        RECT 1234.800 1675.510 1234.940 1685.050 ;
        RECT 1124.340 1675.190 1124.600 1675.510 ;
        RECT 1234.740 1675.190 1235.000 1675.510 ;
        RECT 1124.400 16.730 1124.540 1675.190 ;
        RECT 1120.720 16.590 1124.540 16.730 ;
        RECT 1120.720 2.400 1120.860 16.590 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1145.010 1654.340 1145.330 1654.400 ;
        RECT 1266.450 1654.340 1266.770 1654.400 ;
        RECT 1145.010 1654.200 1266.770 1654.340 ;
        RECT 1145.010 1654.140 1145.330 1654.200 ;
        RECT 1266.450 1654.140 1266.770 1654.200 ;
        RECT 1138.570 19.280 1138.890 19.340 ;
        RECT 1145.010 19.280 1145.330 19.340 ;
        RECT 1138.570 19.140 1145.330 19.280 ;
        RECT 1138.570 19.080 1138.890 19.140 ;
        RECT 1145.010 19.080 1145.330 19.140 ;
      LAYER via ;
        RECT 1145.040 1654.140 1145.300 1654.400 ;
        RECT 1266.480 1654.140 1266.740 1654.400 ;
        RECT 1138.600 19.080 1138.860 19.340 ;
        RECT 1145.040 19.080 1145.300 19.340 ;
      LAYER met2 ;
        RECT 1266.840 1700.410 1267.120 1704.000 ;
        RECT 1266.540 1700.270 1267.120 1700.410 ;
        RECT 1266.540 1654.430 1266.680 1700.270 ;
        RECT 1266.840 1700.000 1267.120 1700.270 ;
        RECT 1145.040 1654.110 1145.300 1654.430 ;
        RECT 1266.480 1654.110 1266.740 1654.430 ;
        RECT 1145.100 19.370 1145.240 1654.110 ;
        RECT 1138.600 19.050 1138.860 19.370 ;
        RECT 1145.040 19.050 1145.300 19.370 ;
        RECT 1138.660 2.400 1138.800 19.050 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1256.330 1684.260 1256.650 1684.320 ;
        RECT 1268.750 1684.260 1269.070 1684.320 ;
        RECT 1256.330 1684.120 1269.070 1684.260 ;
        RECT 1256.330 1684.060 1256.650 1684.120 ;
        RECT 1268.750 1684.060 1269.070 1684.120 ;
        RECT 1156.510 51.580 1156.830 51.640 ;
        RECT 1255.870 51.580 1256.190 51.640 ;
        RECT 1156.510 51.440 1256.190 51.580 ;
        RECT 1156.510 51.380 1156.830 51.440 ;
        RECT 1255.870 51.380 1256.190 51.440 ;
      LAYER via ;
        RECT 1256.360 1684.060 1256.620 1684.320 ;
        RECT 1268.780 1684.060 1269.040 1684.320 ;
        RECT 1156.540 51.380 1156.800 51.640 ;
        RECT 1255.900 51.380 1256.160 51.640 ;
      LAYER met2 ;
        RECT 1268.680 1700.340 1268.960 1704.000 ;
        RECT 1268.680 1700.000 1268.980 1700.340 ;
        RECT 1268.840 1684.350 1268.980 1700.000 ;
        RECT 1256.360 1684.030 1256.620 1684.350 ;
        RECT 1268.780 1684.030 1269.040 1684.350 ;
        RECT 1256.420 1677.290 1256.560 1684.030 ;
        RECT 1255.960 1677.150 1256.560 1677.290 ;
        RECT 1255.960 51.670 1256.100 1677.150 ;
        RECT 1156.540 51.350 1156.800 51.670 ;
        RECT 1255.900 51.350 1256.160 51.670 ;
        RECT 1156.600 2.400 1156.740 51.350 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1215.850 1678.480 1216.170 1678.540 ;
        RECT 1219.070 1678.480 1219.390 1678.540 ;
        RECT 1215.850 1678.340 1219.390 1678.480 ;
        RECT 1215.850 1678.280 1216.170 1678.340 ;
        RECT 1219.070 1678.280 1219.390 1678.340 ;
        RECT 674.430 31.520 674.750 31.580 ;
        RECT 1215.850 31.520 1216.170 31.580 ;
        RECT 674.430 31.380 1216.170 31.520 ;
        RECT 674.430 31.320 674.750 31.380 ;
        RECT 1215.850 31.320 1216.170 31.380 ;
      LAYER via ;
        RECT 1215.880 1678.280 1216.140 1678.540 ;
        RECT 1219.100 1678.280 1219.360 1678.540 ;
        RECT 674.460 31.320 674.720 31.580 ;
        RECT 1215.880 31.320 1216.140 31.580 ;
      LAYER met2 ;
        RECT 1219.000 1700.340 1219.280 1704.000 ;
        RECT 1219.000 1700.000 1219.300 1700.340 ;
        RECT 1219.160 1678.570 1219.300 1700.000 ;
        RECT 1215.880 1678.250 1216.140 1678.570 ;
        RECT 1219.100 1678.250 1219.360 1678.570 ;
        RECT 1215.940 31.610 1216.080 1678.250 ;
        RECT 674.460 31.290 674.720 31.610 ;
        RECT 1215.880 31.290 1216.140 31.610 ;
        RECT 674.520 2.400 674.660 31.290 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1270.590 1679.160 1270.910 1679.220 ;
        RECT 1272.430 1679.160 1272.750 1679.220 ;
        RECT 1270.590 1679.020 1272.750 1679.160 ;
        RECT 1270.590 1678.960 1270.910 1679.020 ;
        RECT 1272.430 1678.960 1272.750 1679.020 ;
        RECT 1173.990 30.840 1174.310 30.900 ;
        RECT 1272.430 30.840 1272.750 30.900 ;
        RECT 1173.990 30.700 1272.750 30.840 ;
        RECT 1173.990 30.640 1174.310 30.700 ;
        RECT 1272.430 30.640 1272.750 30.700 ;
      LAYER via ;
        RECT 1270.620 1678.960 1270.880 1679.220 ;
        RECT 1272.460 1678.960 1272.720 1679.220 ;
        RECT 1174.020 30.640 1174.280 30.900 ;
        RECT 1272.460 30.640 1272.720 30.900 ;
      LAYER met2 ;
        RECT 1270.520 1700.340 1270.800 1704.000 ;
        RECT 1270.520 1700.000 1270.820 1700.340 ;
        RECT 1270.680 1679.250 1270.820 1700.000 ;
        RECT 1270.620 1678.930 1270.880 1679.250 ;
        RECT 1272.460 1678.930 1272.720 1679.250 ;
        RECT 1272.520 30.930 1272.660 1678.930 ;
        RECT 1174.020 30.610 1174.280 30.930 ;
        RECT 1272.460 30.610 1272.720 30.930 ;
        RECT 1174.080 2.400 1174.220 30.610 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1191.930 30.160 1192.250 30.220 ;
        RECT 1271.970 30.160 1272.290 30.220 ;
        RECT 1191.930 30.020 1272.290 30.160 ;
        RECT 1191.930 29.960 1192.250 30.020 ;
        RECT 1271.970 29.960 1272.290 30.020 ;
      LAYER via ;
        RECT 1191.960 29.960 1192.220 30.220 ;
        RECT 1272.000 29.960 1272.260 30.220 ;
      LAYER met2 ;
        RECT 1272.360 1700.410 1272.640 1704.000 ;
        RECT 1272.060 1700.270 1272.640 1700.410 ;
        RECT 1272.060 30.250 1272.200 1700.270 ;
        RECT 1272.360 1700.000 1272.640 1700.270 ;
        RECT 1191.960 29.930 1192.220 30.250 ;
        RECT 1272.000 29.930 1272.260 30.250 ;
        RECT 1192.020 2.400 1192.160 29.930 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1259.090 1645.160 1259.410 1645.220 ;
        RECT 1274.270 1645.160 1274.590 1645.220 ;
        RECT 1259.090 1645.020 1274.590 1645.160 ;
        RECT 1259.090 1644.960 1259.410 1645.020 ;
        RECT 1274.270 1644.960 1274.590 1645.020 ;
        RECT 1209.870 44.780 1210.190 44.840 ;
        RECT 1259.090 44.780 1259.410 44.840 ;
        RECT 1209.870 44.640 1259.410 44.780 ;
        RECT 1209.870 44.580 1210.190 44.640 ;
        RECT 1259.090 44.580 1259.410 44.640 ;
      LAYER via ;
        RECT 1259.120 1644.960 1259.380 1645.220 ;
        RECT 1274.300 1644.960 1274.560 1645.220 ;
        RECT 1209.900 44.580 1210.160 44.840 ;
        RECT 1259.120 44.580 1259.380 44.840 ;
      LAYER met2 ;
        RECT 1274.200 1700.340 1274.480 1704.000 ;
        RECT 1274.200 1700.000 1274.500 1700.340 ;
        RECT 1274.360 1645.250 1274.500 1700.000 ;
        RECT 1259.120 1644.930 1259.380 1645.250 ;
        RECT 1274.300 1644.930 1274.560 1645.250 ;
        RECT 1259.180 44.870 1259.320 1644.930 ;
        RECT 1209.900 44.550 1210.160 44.870 ;
        RECT 1259.120 44.550 1259.380 44.870 ;
        RECT 1209.960 2.400 1210.100 44.550 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 17.920 1228.130 17.980 ;
        RECT 1276.110 17.920 1276.430 17.980 ;
        RECT 1227.810 17.780 1276.430 17.920 ;
        RECT 1227.810 17.720 1228.130 17.780 ;
        RECT 1276.110 17.720 1276.430 17.780 ;
      LAYER via ;
        RECT 1227.840 17.720 1228.100 17.980 ;
        RECT 1276.140 17.720 1276.400 17.980 ;
      LAYER met2 ;
        RECT 1276.040 1700.340 1276.320 1704.000 ;
        RECT 1276.040 1700.000 1276.340 1700.340 ;
        RECT 1276.200 18.010 1276.340 1700.000 ;
        RECT 1227.840 17.690 1228.100 18.010 ;
        RECT 1276.140 17.690 1276.400 18.010 ;
        RECT 1227.900 2.400 1228.040 17.690 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1245.750 14.860 1246.070 14.920 ;
        RECT 1278.410 14.860 1278.730 14.920 ;
        RECT 1245.750 14.720 1278.730 14.860 ;
        RECT 1245.750 14.660 1246.070 14.720 ;
        RECT 1278.410 14.660 1278.730 14.720 ;
      LAYER via ;
        RECT 1245.780 14.660 1246.040 14.920 ;
        RECT 1278.440 14.660 1278.700 14.920 ;
      LAYER met2 ;
        RECT 1277.880 1700.340 1278.160 1704.000 ;
        RECT 1277.880 1700.000 1278.180 1700.340 ;
        RECT 1278.040 1676.610 1278.180 1700.000 ;
        RECT 1278.040 1676.470 1278.640 1676.610 ;
        RECT 1278.500 14.950 1278.640 1676.470 ;
        RECT 1245.780 14.630 1246.040 14.950 ;
        RECT 1278.440 14.630 1278.700 14.950 ;
        RECT 1245.840 2.400 1245.980 14.630 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1279.330 1677.600 1279.650 1677.860 ;
        RECT 1277.490 1675.420 1277.810 1675.480 ;
        RECT 1279.420 1675.420 1279.560 1677.600 ;
        RECT 1277.490 1675.280 1279.560 1675.420 ;
        RECT 1277.490 1675.220 1277.810 1675.280 ;
        RECT 1263.230 17.240 1263.550 17.300 ;
        RECT 1277.490 17.240 1277.810 17.300 ;
        RECT 1263.230 17.100 1277.810 17.240 ;
        RECT 1263.230 17.040 1263.550 17.100 ;
        RECT 1277.490 17.040 1277.810 17.100 ;
      LAYER via ;
        RECT 1279.360 1677.600 1279.620 1677.860 ;
        RECT 1277.520 1675.220 1277.780 1675.480 ;
        RECT 1263.260 17.040 1263.520 17.300 ;
        RECT 1277.520 17.040 1277.780 17.300 ;
      LAYER met2 ;
        RECT 1279.720 1700.410 1280.000 1704.000 ;
        RECT 1279.420 1700.270 1280.000 1700.410 ;
        RECT 1279.420 1677.890 1279.560 1700.270 ;
        RECT 1279.720 1700.000 1280.000 1700.270 ;
        RECT 1279.360 1677.570 1279.620 1677.890 ;
        RECT 1277.520 1675.190 1277.780 1675.510 ;
        RECT 1277.580 17.330 1277.720 1675.190 ;
        RECT 1263.260 17.010 1263.520 17.330 ;
        RECT 1277.520 17.010 1277.780 17.330 ;
        RECT 1263.320 2.400 1263.460 17.010 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.560 1700.340 1281.840 1704.000 ;
        RECT 1281.560 1700.000 1281.860 1700.340 ;
        RECT 1281.720 3.130 1281.860 1700.000 ;
        RECT 1281.260 2.990 1281.860 3.130 ;
        RECT 1281.260 2.400 1281.400 2.990 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1283.470 1685.280 1283.790 1685.340 ;
        RECT 1292.670 1685.280 1292.990 1685.340 ;
        RECT 1283.470 1685.140 1292.990 1685.280 ;
        RECT 1283.470 1685.080 1283.790 1685.140 ;
        RECT 1292.670 1685.080 1292.990 1685.140 ;
        RECT 1292.670 20.640 1292.990 20.700 ;
        RECT 1299.110 20.640 1299.430 20.700 ;
        RECT 1292.670 20.500 1299.430 20.640 ;
        RECT 1292.670 20.440 1292.990 20.500 ;
        RECT 1299.110 20.440 1299.430 20.500 ;
      LAYER via ;
        RECT 1283.500 1685.080 1283.760 1685.340 ;
        RECT 1292.700 1685.080 1292.960 1685.340 ;
        RECT 1292.700 20.440 1292.960 20.700 ;
        RECT 1299.140 20.440 1299.400 20.700 ;
      LAYER met2 ;
        RECT 1283.400 1700.340 1283.680 1704.000 ;
        RECT 1283.400 1700.000 1283.700 1700.340 ;
        RECT 1283.560 1685.370 1283.700 1700.000 ;
        RECT 1283.500 1685.050 1283.760 1685.370 ;
        RECT 1292.700 1685.050 1292.960 1685.370 ;
        RECT 1292.760 20.730 1292.900 1685.050 ;
        RECT 1292.700 20.410 1292.960 20.730 ;
        RECT 1299.140 20.410 1299.400 20.730 ;
        RECT 1299.200 2.400 1299.340 20.410 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1285.310 19.280 1285.630 19.340 ;
        RECT 1317.050 19.280 1317.370 19.340 ;
        RECT 1285.310 19.140 1317.370 19.280 ;
        RECT 1285.310 19.080 1285.630 19.140 ;
        RECT 1317.050 19.080 1317.370 19.140 ;
      LAYER via ;
        RECT 1285.340 19.080 1285.600 19.340 ;
        RECT 1317.080 19.080 1317.340 19.340 ;
      LAYER met2 ;
        RECT 1285.240 1700.340 1285.520 1704.000 ;
        RECT 1285.240 1700.000 1285.540 1700.340 ;
        RECT 1285.400 19.370 1285.540 1700.000 ;
        RECT 1285.340 19.050 1285.600 19.370 ;
        RECT 1317.080 19.050 1317.340 19.370 ;
        RECT 1317.140 2.400 1317.280 19.050 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1287.150 1685.620 1287.470 1685.680 ;
        RECT 1287.150 1685.480 1298.420 1685.620 ;
        RECT 1287.150 1685.420 1287.470 1685.480 ;
        RECT 1298.280 1684.260 1298.420 1685.480 ;
        RECT 1298.280 1684.120 1304.860 1684.260 ;
        RECT 1304.720 1683.240 1304.860 1684.120 ;
        RECT 1305.090 1683.240 1305.410 1683.300 ;
        RECT 1304.720 1683.100 1305.410 1683.240 ;
        RECT 1305.090 1683.040 1305.410 1683.100 ;
        RECT 1305.090 1667.940 1305.410 1668.000 ;
        RECT 1307.850 1667.940 1308.170 1668.000 ;
        RECT 1305.090 1667.800 1308.170 1667.940 ;
        RECT 1305.090 1667.740 1305.410 1667.800 ;
        RECT 1307.850 1667.740 1308.170 1667.800 ;
        RECT 1307.390 41.380 1307.710 41.440 ;
        RECT 1334.990 41.380 1335.310 41.440 ;
        RECT 1307.390 41.240 1335.310 41.380 ;
        RECT 1307.390 41.180 1307.710 41.240 ;
        RECT 1334.990 41.180 1335.310 41.240 ;
      LAYER via ;
        RECT 1287.180 1685.420 1287.440 1685.680 ;
        RECT 1305.120 1683.040 1305.380 1683.300 ;
        RECT 1305.120 1667.740 1305.380 1668.000 ;
        RECT 1307.880 1667.740 1308.140 1668.000 ;
        RECT 1307.420 41.180 1307.680 41.440 ;
        RECT 1335.020 41.180 1335.280 41.440 ;
      LAYER met2 ;
        RECT 1287.080 1700.340 1287.360 1704.000 ;
        RECT 1287.080 1700.000 1287.380 1700.340 ;
        RECT 1287.240 1685.710 1287.380 1700.000 ;
        RECT 1287.180 1685.390 1287.440 1685.710 ;
        RECT 1305.120 1683.010 1305.380 1683.330 ;
        RECT 1305.180 1668.030 1305.320 1683.010 ;
        RECT 1305.120 1667.710 1305.380 1668.030 ;
        RECT 1307.880 1667.710 1308.140 1668.030 ;
        RECT 1307.940 1631.730 1308.080 1667.710 ;
        RECT 1307.480 1631.590 1308.080 1631.730 ;
        RECT 1307.480 41.470 1307.620 1631.590 ;
        RECT 1307.420 41.150 1307.680 41.470 ;
        RECT 1335.020 41.150 1335.280 41.470 ;
        RECT 1335.080 2.400 1335.220 41.150 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 696.510 1639.380 696.830 1639.440 ;
        RECT 1220.910 1639.380 1221.230 1639.440 ;
        RECT 696.510 1639.240 1221.230 1639.380 ;
        RECT 696.510 1639.180 696.830 1639.240 ;
        RECT 1220.910 1639.180 1221.230 1639.240 ;
      LAYER via ;
        RECT 696.540 1639.180 696.800 1639.440 ;
        RECT 1220.940 1639.180 1221.200 1639.440 ;
      LAYER met2 ;
        RECT 1220.840 1700.340 1221.120 1704.000 ;
        RECT 1220.840 1700.000 1221.140 1700.340 ;
        RECT 1221.000 1639.470 1221.140 1700.000 ;
        RECT 696.540 1639.150 696.800 1639.470 ;
        RECT 1220.940 1639.150 1221.200 1639.470 ;
        RECT 696.600 24.210 696.740 1639.150 ;
        RECT 692.460 24.070 696.740 24.210 ;
        RECT 692.460 2.400 692.600 24.070 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1288.990 27.440 1289.310 27.500 ;
        RECT 1352.930 27.440 1353.250 27.500 ;
        RECT 1288.990 27.300 1353.250 27.440 ;
        RECT 1288.990 27.240 1289.310 27.300 ;
        RECT 1352.930 27.240 1353.250 27.300 ;
      LAYER via ;
        RECT 1289.020 27.240 1289.280 27.500 ;
        RECT 1352.960 27.240 1353.220 27.500 ;
      LAYER met2 ;
        RECT 1288.920 1700.340 1289.200 1704.000 ;
        RECT 1288.920 1700.000 1289.220 1700.340 ;
        RECT 1289.080 27.530 1289.220 1700.000 ;
        RECT 1289.020 27.210 1289.280 27.530 ;
        RECT 1352.960 27.210 1353.220 27.530 ;
        RECT 1353.020 5.170 1353.160 27.210 ;
        RECT 1352.560 5.030 1353.160 5.170 ;
        RECT 1352.560 2.400 1352.700 5.030 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1290.830 1683.920 1291.150 1683.980 ;
        RECT 1293.130 1683.920 1293.450 1683.980 ;
        RECT 1290.830 1683.780 1293.450 1683.920 ;
        RECT 1290.830 1683.720 1291.150 1683.780 ;
        RECT 1293.130 1683.720 1293.450 1683.780 ;
        RECT 1293.130 27.100 1293.450 27.160 ;
        RECT 1370.410 27.100 1370.730 27.160 ;
        RECT 1293.130 26.960 1370.730 27.100 ;
        RECT 1293.130 26.900 1293.450 26.960 ;
        RECT 1370.410 26.900 1370.730 26.960 ;
      LAYER via ;
        RECT 1290.860 1683.720 1291.120 1683.980 ;
        RECT 1293.160 1683.720 1293.420 1683.980 ;
        RECT 1293.160 26.900 1293.420 27.160 ;
        RECT 1370.440 26.900 1370.700 27.160 ;
      LAYER met2 ;
        RECT 1290.760 1700.340 1291.040 1704.000 ;
        RECT 1290.760 1700.000 1291.060 1700.340 ;
        RECT 1290.920 1684.010 1291.060 1700.000 ;
        RECT 1290.860 1683.690 1291.120 1684.010 ;
        RECT 1293.160 1683.690 1293.420 1684.010 ;
        RECT 1293.220 27.190 1293.360 1683.690 ;
        RECT 1293.160 26.870 1293.420 27.190 ;
        RECT 1370.440 26.870 1370.700 27.190 ;
        RECT 1370.500 2.400 1370.640 26.870 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1292.210 26.080 1292.530 26.140 ;
        RECT 1388.350 26.080 1388.670 26.140 ;
        RECT 1292.210 25.940 1388.670 26.080 ;
        RECT 1292.210 25.880 1292.530 25.940 ;
        RECT 1388.350 25.880 1388.670 25.940 ;
      LAYER via ;
        RECT 1292.240 25.880 1292.500 26.140 ;
        RECT 1388.380 25.880 1388.640 26.140 ;
      LAYER met2 ;
        RECT 1292.600 1700.410 1292.880 1704.000 ;
        RECT 1292.300 1700.270 1292.880 1700.410 ;
        RECT 1292.300 26.170 1292.440 1700.270 ;
        RECT 1292.600 1700.000 1292.880 1700.270 ;
        RECT 1292.240 25.850 1292.500 26.170 ;
        RECT 1388.380 25.850 1388.640 26.170 ;
        RECT 1388.440 2.400 1388.580 25.850 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1294.510 1684.260 1294.830 1684.320 ;
        RECT 1296.350 1684.260 1296.670 1684.320 ;
        RECT 1294.510 1684.120 1296.670 1684.260 ;
        RECT 1294.510 1684.060 1294.830 1684.120 ;
        RECT 1296.350 1684.060 1296.670 1684.120 ;
        RECT 1296.350 25.400 1296.670 25.460 ;
        RECT 1406.290 25.400 1406.610 25.460 ;
        RECT 1296.350 25.260 1406.610 25.400 ;
        RECT 1296.350 25.200 1296.670 25.260 ;
        RECT 1406.290 25.200 1406.610 25.260 ;
      LAYER via ;
        RECT 1294.540 1684.060 1294.800 1684.320 ;
        RECT 1296.380 1684.060 1296.640 1684.320 ;
        RECT 1296.380 25.200 1296.640 25.460 ;
        RECT 1406.320 25.200 1406.580 25.460 ;
      LAYER met2 ;
        RECT 1294.440 1700.340 1294.720 1704.000 ;
        RECT 1294.440 1700.000 1294.740 1700.340 ;
        RECT 1294.600 1684.350 1294.740 1700.000 ;
        RECT 1294.540 1684.030 1294.800 1684.350 ;
        RECT 1296.380 1684.030 1296.640 1684.350 ;
        RECT 1296.440 25.490 1296.580 1684.030 ;
        RECT 1296.380 25.170 1296.640 25.490 ;
        RECT 1406.320 25.170 1406.580 25.490 ;
        RECT 1406.380 2.400 1406.520 25.170 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1295.890 25.060 1296.210 25.120 ;
        RECT 1423.770 25.060 1424.090 25.120 ;
        RECT 1295.890 24.920 1424.090 25.060 ;
        RECT 1295.890 24.860 1296.210 24.920 ;
        RECT 1423.770 24.860 1424.090 24.920 ;
      LAYER via ;
        RECT 1295.920 24.860 1296.180 25.120 ;
        RECT 1423.800 24.860 1424.060 25.120 ;
      LAYER met2 ;
        RECT 1296.280 1700.410 1296.560 1704.000 ;
        RECT 1295.980 1700.270 1296.560 1700.410 ;
        RECT 1295.980 25.150 1296.120 1700.270 ;
        RECT 1296.280 1700.000 1296.560 1700.270 ;
        RECT 1295.920 24.830 1296.180 25.150 ;
        RECT 1423.800 24.830 1424.060 25.150 ;
        RECT 1423.860 2.400 1424.000 24.830 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1298.190 1686.300 1298.510 1686.360 ;
        RECT 1311.070 1686.300 1311.390 1686.360 ;
        RECT 1298.190 1686.160 1311.390 1686.300 ;
        RECT 1298.190 1686.100 1298.510 1686.160 ;
        RECT 1311.070 1686.100 1311.390 1686.160 ;
        RECT 1311.070 1673.040 1311.390 1673.100 ;
        RECT 1435.270 1673.040 1435.590 1673.100 ;
        RECT 1311.070 1672.900 1435.590 1673.040 ;
        RECT 1311.070 1672.840 1311.390 1672.900 ;
        RECT 1435.270 1672.840 1435.590 1672.900 ;
        RECT 1435.270 20.980 1435.590 21.040 ;
        RECT 1441.710 20.980 1442.030 21.040 ;
        RECT 1435.270 20.840 1442.030 20.980 ;
        RECT 1435.270 20.780 1435.590 20.840 ;
        RECT 1441.710 20.780 1442.030 20.840 ;
      LAYER via ;
        RECT 1298.220 1686.100 1298.480 1686.360 ;
        RECT 1311.100 1686.100 1311.360 1686.360 ;
        RECT 1311.100 1672.840 1311.360 1673.100 ;
        RECT 1435.300 1672.840 1435.560 1673.100 ;
        RECT 1435.300 20.780 1435.560 21.040 ;
        RECT 1441.740 20.780 1442.000 21.040 ;
      LAYER met2 ;
        RECT 1298.120 1700.340 1298.400 1704.000 ;
        RECT 1298.120 1700.000 1298.420 1700.340 ;
        RECT 1298.280 1686.390 1298.420 1700.000 ;
        RECT 1298.220 1686.070 1298.480 1686.390 ;
        RECT 1311.100 1686.070 1311.360 1686.390 ;
        RECT 1311.160 1673.130 1311.300 1686.070 ;
        RECT 1311.100 1672.810 1311.360 1673.130 ;
        RECT 1435.300 1672.810 1435.560 1673.130 ;
        RECT 1435.360 21.070 1435.500 1672.810 ;
        RECT 1435.300 20.750 1435.560 21.070 ;
        RECT 1441.740 20.750 1442.000 21.070 ;
        RECT 1441.800 2.400 1441.940 20.750 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1299.645 1228.165 1299.815 1276.275 ;
        RECT 1299.645 462.485 1299.815 476.255 ;
      LAYER mcon ;
        RECT 1299.645 1276.105 1299.815 1276.275 ;
        RECT 1299.645 476.085 1299.815 476.255 ;
      LAYER met1 ;
        RECT 1299.570 1353.100 1299.890 1353.160 ;
        RECT 1299.200 1352.960 1299.890 1353.100 ;
        RECT 1299.200 1352.480 1299.340 1352.960 ;
        RECT 1299.570 1352.900 1299.890 1352.960 ;
        RECT 1299.110 1352.220 1299.430 1352.480 ;
        RECT 1299.570 1276.260 1299.890 1276.320 ;
        RECT 1299.375 1276.120 1299.890 1276.260 ;
        RECT 1299.570 1276.060 1299.890 1276.120 ;
        RECT 1299.570 1228.320 1299.890 1228.380 ;
        RECT 1299.375 1228.180 1299.890 1228.320 ;
        RECT 1299.570 1228.120 1299.890 1228.180 ;
        RECT 1299.110 1028.200 1299.430 1028.460 ;
        RECT 1299.200 1028.060 1299.340 1028.200 ;
        RECT 1299.570 1028.060 1299.890 1028.120 ;
        RECT 1299.200 1027.920 1299.890 1028.060 ;
        RECT 1299.570 1027.860 1299.890 1027.920 ;
        RECT 1299.570 848.880 1299.890 848.940 ;
        RECT 1298.740 848.740 1299.890 848.880 ;
        RECT 1298.740 848.600 1298.880 848.740 ;
        RECT 1299.570 848.680 1299.890 848.740 ;
        RECT 1298.650 848.340 1298.970 848.600 ;
        RECT 1298.650 800.600 1298.970 800.660 ;
        RECT 1299.570 800.600 1299.890 800.660 ;
        RECT 1298.650 800.460 1299.890 800.600 ;
        RECT 1298.650 800.400 1298.970 800.460 ;
        RECT 1299.570 800.400 1299.890 800.460 ;
        RECT 1299.110 738.180 1299.430 738.440 ;
        RECT 1299.200 738.040 1299.340 738.180 ;
        RECT 1299.570 738.040 1299.890 738.100 ;
        RECT 1299.200 737.900 1299.890 738.040 ;
        RECT 1299.570 737.840 1299.890 737.900 ;
        RECT 1299.110 641.620 1299.430 641.880 ;
        RECT 1299.200 641.480 1299.340 641.620 ;
        RECT 1299.570 641.480 1299.890 641.540 ;
        RECT 1299.200 641.340 1299.890 641.480 ;
        RECT 1299.570 641.280 1299.890 641.340 ;
        RECT 1299.110 579.600 1299.430 579.660 ;
        RECT 1299.570 579.600 1299.890 579.660 ;
        RECT 1299.110 579.460 1299.890 579.600 ;
        RECT 1299.110 579.400 1299.430 579.460 ;
        RECT 1299.570 579.400 1299.890 579.460 ;
        RECT 1299.570 476.240 1299.890 476.300 ;
        RECT 1299.375 476.100 1299.890 476.240 ;
        RECT 1299.570 476.040 1299.890 476.100 ;
        RECT 1299.570 462.640 1299.890 462.700 ;
        RECT 1299.375 462.500 1299.890 462.640 ;
        RECT 1299.570 462.440 1299.890 462.500 ;
        RECT 1299.110 407.220 1299.430 407.280 ;
        RECT 1299.570 407.220 1299.890 407.280 ;
        RECT 1299.110 407.080 1299.890 407.220 ;
        RECT 1299.110 407.020 1299.430 407.080 ;
        RECT 1299.570 407.020 1299.890 407.080 ;
        RECT 1299.110 365.740 1299.430 365.800 ;
        RECT 1300.490 365.740 1300.810 365.800 ;
        RECT 1299.110 365.600 1300.810 365.740 ;
        RECT 1299.110 365.540 1299.430 365.600 ;
        RECT 1300.490 365.540 1300.810 365.600 ;
        RECT 1298.650 310.660 1298.970 310.720 ;
        RECT 1299.110 310.660 1299.430 310.720 ;
        RECT 1298.650 310.520 1299.430 310.660 ;
        RECT 1298.650 310.460 1298.970 310.520 ;
        RECT 1299.110 310.460 1299.430 310.520 ;
        RECT 1299.110 255.380 1299.430 255.640 ;
        RECT 1299.200 255.240 1299.340 255.380 ;
        RECT 1299.570 255.240 1299.890 255.300 ;
        RECT 1299.200 255.100 1299.890 255.240 ;
        RECT 1299.570 255.040 1299.890 255.100 ;
        RECT 1299.110 137.940 1299.430 138.000 ;
        RECT 1299.570 137.940 1299.890 138.000 ;
        RECT 1299.110 137.800 1299.890 137.940 ;
        RECT 1299.110 137.740 1299.430 137.800 ;
        RECT 1299.570 137.740 1299.890 137.800 ;
        RECT 1299.570 46.480 1299.890 46.540 ;
        RECT 1459.650 46.480 1459.970 46.540 ;
        RECT 1299.570 46.340 1459.970 46.480 ;
        RECT 1299.570 46.280 1299.890 46.340 ;
        RECT 1459.650 46.280 1459.970 46.340 ;
      LAYER via ;
        RECT 1299.600 1352.900 1299.860 1353.160 ;
        RECT 1299.140 1352.220 1299.400 1352.480 ;
        RECT 1299.600 1276.060 1299.860 1276.320 ;
        RECT 1299.600 1228.120 1299.860 1228.380 ;
        RECT 1299.140 1028.200 1299.400 1028.460 ;
        RECT 1299.600 1027.860 1299.860 1028.120 ;
        RECT 1299.600 848.680 1299.860 848.940 ;
        RECT 1298.680 848.340 1298.940 848.600 ;
        RECT 1298.680 800.400 1298.940 800.660 ;
        RECT 1299.600 800.400 1299.860 800.660 ;
        RECT 1299.140 738.180 1299.400 738.440 ;
        RECT 1299.600 737.840 1299.860 738.100 ;
        RECT 1299.140 641.620 1299.400 641.880 ;
        RECT 1299.600 641.280 1299.860 641.540 ;
        RECT 1299.140 579.400 1299.400 579.660 ;
        RECT 1299.600 579.400 1299.860 579.660 ;
        RECT 1299.600 476.040 1299.860 476.300 ;
        RECT 1299.600 462.440 1299.860 462.700 ;
        RECT 1299.140 407.020 1299.400 407.280 ;
        RECT 1299.600 407.020 1299.860 407.280 ;
        RECT 1299.140 365.540 1299.400 365.800 ;
        RECT 1300.520 365.540 1300.780 365.800 ;
        RECT 1298.680 310.460 1298.940 310.720 ;
        RECT 1299.140 310.460 1299.400 310.720 ;
        RECT 1299.140 255.380 1299.400 255.640 ;
        RECT 1299.600 255.040 1299.860 255.300 ;
        RECT 1299.140 137.740 1299.400 138.000 ;
        RECT 1299.600 137.740 1299.860 138.000 ;
        RECT 1299.600 46.280 1299.860 46.540 ;
        RECT 1459.680 46.280 1459.940 46.540 ;
      LAYER met2 ;
        RECT 1299.960 1700.410 1300.240 1704.000 ;
        RECT 1299.660 1700.270 1300.240 1700.410 ;
        RECT 1299.660 1659.610 1299.800 1700.270 ;
        RECT 1299.960 1700.000 1300.240 1700.270 ;
        RECT 1299.200 1659.470 1299.800 1659.610 ;
        RECT 1299.200 1507.970 1299.340 1659.470 ;
        RECT 1299.200 1507.830 1299.800 1507.970 ;
        RECT 1299.660 1353.190 1299.800 1507.830 ;
        RECT 1299.600 1352.870 1299.860 1353.190 ;
        RECT 1299.140 1352.190 1299.400 1352.510 ;
        RECT 1299.200 1321.650 1299.340 1352.190 ;
        RECT 1299.200 1321.510 1299.800 1321.650 ;
        RECT 1299.660 1276.350 1299.800 1321.510 ;
        RECT 1299.600 1276.030 1299.860 1276.350 ;
        RECT 1299.600 1228.090 1299.860 1228.410 ;
        RECT 1299.660 1087.050 1299.800 1228.090 ;
        RECT 1299.200 1086.910 1299.800 1087.050 ;
        RECT 1299.200 1028.490 1299.340 1086.910 ;
        RECT 1299.140 1028.170 1299.400 1028.490 ;
        RECT 1299.600 1027.830 1299.860 1028.150 ;
        RECT 1299.660 945.725 1299.800 1027.830 ;
        RECT 1299.590 945.355 1299.870 945.725 ;
        RECT 1298.670 944.930 1298.950 945.045 ;
        RECT 1298.670 944.790 1299.340 944.930 ;
        RECT 1298.670 944.675 1298.950 944.790 ;
        RECT 1299.200 910.250 1299.340 944.790 ;
        RECT 1299.200 910.110 1299.800 910.250 ;
        RECT 1299.660 848.970 1299.800 910.110 ;
        RECT 1299.600 848.650 1299.860 848.970 ;
        RECT 1298.680 848.310 1298.940 848.630 ;
        RECT 1298.740 800.690 1298.880 848.310 ;
        RECT 1298.680 800.370 1298.940 800.690 ;
        RECT 1299.600 800.370 1299.860 800.690 ;
        RECT 1299.660 787.170 1299.800 800.370 ;
        RECT 1299.200 787.030 1299.800 787.170 ;
        RECT 1299.200 738.470 1299.340 787.030 ;
        RECT 1299.140 738.150 1299.400 738.470 ;
        RECT 1299.600 737.810 1299.860 738.130 ;
        RECT 1299.660 690.610 1299.800 737.810 ;
        RECT 1299.200 690.470 1299.800 690.610 ;
        RECT 1299.200 641.910 1299.340 690.470 ;
        RECT 1299.140 641.590 1299.400 641.910 ;
        RECT 1299.600 641.250 1299.860 641.570 ;
        RECT 1299.660 603.570 1299.800 641.250 ;
        RECT 1299.200 603.430 1299.800 603.570 ;
        RECT 1299.200 579.690 1299.340 603.430 ;
        RECT 1299.140 579.370 1299.400 579.690 ;
        RECT 1299.600 579.370 1299.860 579.690 ;
        RECT 1299.660 476.330 1299.800 579.370 ;
        RECT 1299.600 476.010 1299.860 476.330 ;
        RECT 1299.600 462.410 1299.860 462.730 ;
        RECT 1299.660 407.310 1299.800 462.410 ;
        RECT 1299.140 406.990 1299.400 407.310 ;
        RECT 1299.600 406.990 1299.860 407.310 ;
        RECT 1299.200 365.830 1299.340 406.990 ;
        RECT 1299.140 365.510 1299.400 365.830 ;
        RECT 1300.520 365.510 1300.780 365.830 ;
        RECT 1300.580 358.885 1300.720 365.510 ;
        RECT 1298.670 358.515 1298.950 358.885 ;
        RECT 1300.510 358.515 1300.790 358.885 ;
        RECT 1298.740 310.750 1298.880 358.515 ;
        RECT 1298.680 310.430 1298.940 310.750 ;
        RECT 1299.140 310.430 1299.400 310.750 ;
        RECT 1299.200 255.670 1299.340 310.430 ;
        RECT 1299.140 255.350 1299.400 255.670 ;
        RECT 1299.600 255.010 1299.860 255.330 ;
        RECT 1299.660 217.330 1299.800 255.010 ;
        RECT 1299.200 217.190 1299.800 217.330 ;
        RECT 1299.200 138.030 1299.340 217.190 ;
        RECT 1299.140 137.710 1299.400 138.030 ;
        RECT 1299.600 137.710 1299.860 138.030 ;
        RECT 1299.660 46.570 1299.800 137.710 ;
        RECT 1299.600 46.250 1299.860 46.570 ;
        RECT 1459.680 46.250 1459.940 46.570 ;
        RECT 1459.740 2.400 1459.880 46.250 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
      LAYER via2 ;
        RECT 1299.590 945.400 1299.870 945.680 ;
        RECT 1298.670 944.720 1298.950 945.000 ;
        RECT 1298.670 358.560 1298.950 358.840 ;
        RECT 1300.510 358.560 1300.790 358.840 ;
      LAYER met3 ;
        RECT 1299.565 945.690 1299.895 945.705 ;
        RECT 1298.660 945.390 1299.895 945.690 ;
        RECT 1298.660 945.025 1298.960 945.390 ;
        RECT 1299.565 945.375 1299.895 945.390 ;
        RECT 1298.645 944.695 1298.975 945.025 ;
        RECT 1298.645 358.850 1298.975 358.865 ;
        RECT 1300.485 358.850 1300.815 358.865 ;
        RECT 1298.645 358.550 1300.815 358.850 ;
        RECT 1298.645 358.535 1298.975 358.550 ;
        RECT 1300.485 358.535 1300.815 358.550 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1300.030 317.600 1300.350 317.860 ;
        RECT 1300.120 317.180 1300.260 317.600 ;
        RECT 1300.030 316.920 1300.350 317.180 ;
        RECT 1300.030 46.140 1300.350 46.200 ;
        RECT 1477.590 46.140 1477.910 46.200 ;
        RECT 1300.030 46.000 1477.910 46.140 ;
        RECT 1300.030 45.940 1300.350 46.000 ;
        RECT 1477.590 45.940 1477.910 46.000 ;
      LAYER via ;
        RECT 1300.060 317.600 1300.320 317.860 ;
        RECT 1300.060 316.920 1300.320 317.180 ;
        RECT 1300.060 45.940 1300.320 46.200 ;
        RECT 1477.620 45.940 1477.880 46.200 ;
      LAYER met2 ;
        RECT 1301.340 1700.340 1301.620 1704.000 ;
        RECT 1301.340 1700.000 1301.640 1700.340 ;
        RECT 1301.500 1678.140 1301.640 1700.000 ;
        RECT 1300.120 1678.000 1301.640 1678.140 ;
        RECT 1300.120 317.890 1300.260 1678.000 ;
        RECT 1300.060 317.570 1300.320 317.890 ;
        RECT 1300.060 316.890 1300.320 317.210 ;
        RECT 1300.120 46.230 1300.260 316.890 ;
        RECT 1300.060 45.910 1300.320 46.230 ;
        RECT 1477.620 45.910 1477.880 46.230 ;
        RECT 1477.680 2.400 1477.820 45.910 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1303.325 1573.265 1303.495 1609.475 ;
        RECT 1302.865 1187.025 1303.035 1235.135 ;
        RECT 1303.325 938.485 1303.495 985.915 ;
        RECT 1303.325 890.205 1303.495 897.175 ;
        RECT 1302.865 745.365 1303.035 793.475 ;
        RECT 1302.865 648.805 1303.035 703.715 ;
        RECT 1302.405 510.425 1302.575 552.075 ;
        RECT 1303.325 45.645 1303.495 82.875 ;
      LAYER mcon ;
        RECT 1303.325 1609.305 1303.495 1609.475 ;
        RECT 1302.865 1234.965 1303.035 1235.135 ;
        RECT 1303.325 985.745 1303.495 985.915 ;
        RECT 1303.325 897.005 1303.495 897.175 ;
        RECT 1302.865 793.305 1303.035 793.475 ;
        RECT 1302.865 703.545 1303.035 703.715 ;
        RECT 1302.405 551.905 1302.575 552.075 ;
        RECT 1303.325 82.705 1303.495 82.875 ;
      LAYER met1 ;
        RECT 1301.870 1621.700 1302.190 1621.760 ;
        RECT 1303.250 1621.700 1303.570 1621.760 ;
        RECT 1301.870 1621.560 1303.570 1621.700 ;
        RECT 1301.870 1621.500 1302.190 1621.560 ;
        RECT 1303.250 1621.500 1303.570 1621.560 ;
        RECT 1303.250 1609.460 1303.570 1609.520 ;
        RECT 1303.055 1609.320 1303.570 1609.460 ;
        RECT 1303.250 1609.260 1303.570 1609.320 ;
        RECT 1303.250 1573.420 1303.570 1573.480 ;
        RECT 1303.055 1573.280 1303.570 1573.420 ;
        RECT 1303.250 1573.220 1303.570 1573.280 ;
        RECT 1302.805 1235.120 1303.095 1235.165 ;
        RECT 1303.250 1235.120 1303.570 1235.180 ;
        RECT 1302.805 1234.980 1303.570 1235.120 ;
        RECT 1302.805 1234.935 1303.095 1234.980 ;
        RECT 1303.250 1234.920 1303.570 1234.980 ;
        RECT 1302.790 1187.180 1303.110 1187.240 ;
        RECT 1302.595 1187.040 1303.110 1187.180 ;
        RECT 1302.790 1186.980 1303.110 1187.040 ;
        RECT 1303.710 1097.420 1304.030 1097.480 ;
        RECT 1303.340 1097.280 1304.030 1097.420 ;
        RECT 1303.340 1097.140 1303.480 1097.280 ;
        RECT 1303.710 1097.220 1304.030 1097.280 ;
        RECT 1303.250 1096.880 1303.570 1097.140 ;
        RECT 1303.250 1089.940 1303.570 1090.000 ;
        RECT 1304.630 1089.940 1304.950 1090.000 ;
        RECT 1303.250 1089.800 1304.950 1089.940 ;
        RECT 1303.250 1089.740 1303.570 1089.800 ;
        RECT 1304.630 1089.740 1304.950 1089.800 ;
        RECT 1303.250 993.380 1303.570 993.440 ;
        RECT 1303.710 993.380 1304.030 993.440 ;
        RECT 1303.250 993.240 1304.030 993.380 ;
        RECT 1303.250 993.180 1303.570 993.240 ;
        RECT 1303.710 993.180 1304.030 993.240 ;
        RECT 1303.250 986.380 1303.570 986.640 ;
        RECT 1303.340 985.945 1303.480 986.380 ;
        RECT 1303.265 985.715 1303.555 985.945 ;
        RECT 1303.250 938.640 1303.570 938.700 ;
        RECT 1303.055 938.500 1303.570 938.640 ;
        RECT 1303.250 938.440 1303.570 938.500 ;
        RECT 1303.250 897.160 1303.570 897.220 ;
        RECT 1303.055 897.020 1303.570 897.160 ;
        RECT 1303.250 896.960 1303.570 897.020 ;
        RECT 1303.250 890.360 1303.570 890.420 ;
        RECT 1303.055 890.220 1303.570 890.360 ;
        RECT 1303.250 890.160 1303.570 890.220 ;
        RECT 1302.790 793.460 1303.110 793.520 ;
        RECT 1302.595 793.320 1303.110 793.460 ;
        RECT 1302.790 793.260 1303.110 793.320 ;
        RECT 1302.805 745.520 1303.095 745.565 ;
        RECT 1303.250 745.520 1303.570 745.580 ;
        RECT 1302.805 745.380 1303.570 745.520 ;
        RECT 1302.805 745.335 1303.095 745.380 ;
        RECT 1303.250 745.320 1303.570 745.380 ;
        RECT 1302.790 703.700 1303.110 703.760 ;
        RECT 1302.595 703.560 1303.110 703.700 ;
        RECT 1302.790 703.500 1303.110 703.560 ;
        RECT 1302.790 648.960 1303.110 649.020 ;
        RECT 1302.595 648.820 1303.110 648.960 ;
        RECT 1302.790 648.760 1303.110 648.820 ;
        RECT 1302.330 558.860 1302.650 558.920 ;
        RECT 1302.790 558.860 1303.110 558.920 ;
        RECT 1302.330 558.720 1303.110 558.860 ;
        RECT 1302.330 558.660 1302.650 558.720 ;
        RECT 1302.790 558.660 1303.110 558.720 ;
        RECT 1302.330 552.060 1302.650 552.120 ;
        RECT 1302.135 551.920 1302.650 552.060 ;
        RECT 1302.330 551.860 1302.650 551.920 ;
        RECT 1302.345 510.580 1302.635 510.625 ;
        RECT 1302.790 510.580 1303.110 510.640 ;
        RECT 1302.345 510.440 1303.110 510.580 ;
        RECT 1302.345 510.395 1302.635 510.440 ;
        RECT 1302.790 510.380 1303.110 510.440 ;
        RECT 1302.790 227.500 1303.110 227.760 ;
        RECT 1302.880 227.080 1303.020 227.500 ;
        RECT 1302.790 226.820 1303.110 227.080 ;
        RECT 1302.790 173.100 1303.110 173.360 ;
        RECT 1302.880 172.620 1303.020 173.100 ;
        RECT 1303.250 172.620 1303.570 172.680 ;
        RECT 1302.880 172.480 1303.570 172.620 ;
        RECT 1303.250 172.420 1303.570 172.480 ;
        RECT 1303.250 145.080 1303.570 145.140 ;
        RECT 1302.880 144.940 1303.570 145.080 ;
        RECT 1302.880 144.800 1303.020 144.940 ;
        RECT 1303.250 144.880 1303.570 144.940 ;
        RECT 1302.790 144.540 1303.110 144.800 ;
        RECT 1303.250 82.860 1303.570 82.920 ;
        RECT 1303.055 82.720 1303.570 82.860 ;
        RECT 1303.250 82.660 1303.570 82.720 ;
        RECT 1303.265 45.800 1303.555 45.845 ;
        RECT 1495.530 45.800 1495.850 45.860 ;
        RECT 1303.265 45.660 1495.850 45.800 ;
        RECT 1303.265 45.615 1303.555 45.660 ;
        RECT 1495.530 45.600 1495.850 45.660 ;
      LAYER via ;
        RECT 1301.900 1621.500 1302.160 1621.760 ;
        RECT 1303.280 1621.500 1303.540 1621.760 ;
        RECT 1303.280 1609.260 1303.540 1609.520 ;
        RECT 1303.280 1573.220 1303.540 1573.480 ;
        RECT 1303.280 1234.920 1303.540 1235.180 ;
        RECT 1302.820 1186.980 1303.080 1187.240 ;
        RECT 1303.740 1097.220 1304.000 1097.480 ;
        RECT 1303.280 1096.880 1303.540 1097.140 ;
        RECT 1303.280 1089.740 1303.540 1090.000 ;
        RECT 1304.660 1089.740 1304.920 1090.000 ;
        RECT 1303.280 993.180 1303.540 993.440 ;
        RECT 1303.740 993.180 1304.000 993.440 ;
        RECT 1303.280 986.380 1303.540 986.640 ;
        RECT 1303.280 938.440 1303.540 938.700 ;
        RECT 1303.280 896.960 1303.540 897.220 ;
        RECT 1303.280 890.160 1303.540 890.420 ;
        RECT 1302.820 793.260 1303.080 793.520 ;
        RECT 1303.280 745.320 1303.540 745.580 ;
        RECT 1302.820 703.500 1303.080 703.760 ;
        RECT 1302.820 648.760 1303.080 649.020 ;
        RECT 1302.360 558.660 1302.620 558.920 ;
        RECT 1302.820 558.660 1303.080 558.920 ;
        RECT 1302.360 551.860 1302.620 552.120 ;
        RECT 1302.820 510.380 1303.080 510.640 ;
        RECT 1302.820 227.500 1303.080 227.760 ;
        RECT 1302.820 226.820 1303.080 227.080 ;
        RECT 1302.820 173.100 1303.080 173.360 ;
        RECT 1303.280 172.420 1303.540 172.680 ;
        RECT 1303.280 144.880 1303.540 145.140 ;
        RECT 1302.820 144.540 1303.080 144.800 ;
        RECT 1303.280 82.660 1303.540 82.920 ;
        RECT 1495.560 45.600 1495.820 45.860 ;
      LAYER met2 ;
        RECT 1303.180 1700.340 1303.460 1704.000 ;
        RECT 1303.180 1700.000 1303.480 1700.340 ;
        RECT 1303.340 1621.790 1303.480 1700.000 ;
        RECT 1301.900 1621.645 1302.160 1621.790 ;
        RECT 1303.280 1621.645 1303.540 1621.790 ;
        RECT 1301.890 1621.275 1302.170 1621.645 ;
        RECT 1303.270 1621.275 1303.550 1621.645 ;
        RECT 1303.340 1609.550 1303.480 1621.275 ;
        RECT 1303.280 1609.230 1303.540 1609.550 ;
        RECT 1303.280 1573.190 1303.540 1573.510 ;
        RECT 1303.340 1332.645 1303.480 1573.190 ;
        RECT 1303.270 1332.275 1303.550 1332.645 ;
        RECT 1303.270 1331.595 1303.550 1331.965 ;
        RECT 1303.340 1235.210 1303.480 1331.595 ;
        RECT 1303.280 1234.890 1303.540 1235.210 ;
        RECT 1302.820 1186.950 1303.080 1187.270 ;
        RECT 1302.880 1138.845 1303.020 1186.950 ;
        RECT 1302.810 1138.475 1303.090 1138.845 ;
        RECT 1303.730 1138.475 1304.010 1138.845 ;
        RECT 1303.800 1097.510 1303.940 1138.475 ;
        RECT 1303.740 1097.190 1304.000 1097.510 ;
        RECT 1303.280 1096.850 1303.540 1097.170 ;
        RECT 1303.340 1090.030 1303.480 1096.850 ;
        RECT 1303.280 1089.710 1303.540 1090.030 ;
        RECT 1304.660 1089.710 1304.920 1090.030 ;
        RECT 1304.720 1042.285 1304.860 1089.710 ;
        RECT 1304.650 1041.915 1304.930 1042.285 ;
        RECT 1303.730 1041.235 1304.010 1041.605 ;
        RECT 1303.800 993.470 1303.940 1041.235 ;
        RECT 1303.280 993.150 1303.540 993.470 ;
        RECT 1303.740 993.150 1304.000 993.470 ;
        RECT 1303.340 986.670 1303.480 993.150 ;
        RECT 1303.280 986.350 1303.540 986.670 ;
        RECT 1303.280 938.410 1303.540 938.730 ;
        RECT 1303.340 897.250 1303.480 938.410 ;
        RECT 1303.280 896.930 1303.540 897.250 ;
        RECT 1303.280 890.130 1303.540 890.450 ;
        RECT 1303.340 889.965 1303.480 890.130 ;
        RECT 1303.270 889.595 1303.550 889.965 ;
        RECT 1304.190 889.595 1304.470 889.965 ;
        RECT 1304.260 842.365 1304.400 889.595 ;
        RECT 1303.270 841.995 1303.550 842.365 ;
        RECT 1304.190 841.995 1304.470 842.365 ;
        RECT 1303.340 814.370 1303.480 841.995 ;
        RECT 1302.880 814.230 1303.480 814.370 ;
        RECT 1302.880 793.550 1303.020 814.230 ;
        RECT 1302.820 793.230 1303.080 793.550 ;
        RECT 1303.280 745.290 1303.540 745.610 ;
        RECT 1303.340 704.210 1303.480 745.290 ;
        RECT 1302.880 704.070 1303.480 704.210 ;
        RECT 1302.880 703.790 1303.020 704.070 ;
        RECT 1302.820 703.470 1303.080 703.790 ;
        RECT 1302.820 648.730 1303.080 649.050 ;
        RECT 1302.880 558.950 1303.020 648.730 ;
        RECT 1302.360 558.630 1302.620 558.950 ;
        RECT 1302.820 558.630 1303.080 558.950 ;
        RECT 1302.420 552.150 1302.560 558.630 ;
        RECT 1302.360 551.830 1302.620 552.150 ;
        RECT 1302.820 510.350 1303.080 510.670 ;
        RECT 1302.880 503.725 1303.020 510.350 ;
        RECT 1302.810 503.355 1303.090 503.725 ;
        RECT 1303.270 502.675 1303.550 503.045 ;
        RECT 1303.340 390.050 1303.480 502.675 ;
        RECT 1302.880 389.910 1303.480 390.050 ;
        RECT 1302.880 227.790 1303.020 389.910 ;
        RECT 1302.820 227.470 1303.080 227.790 ;
        RECT 1302.820 226.790 1303.080 227.110 ;
        RECT 1302.880 173.390 1303.020 226.790 ;
        RECT 1302.820 173.070 1303.080 173.390 ;
        RECT 1303.280 172.390 1303.540 172.710 ;
        RECT 1303.340 145.170 1303.480 172.390 ;
        RECT 1303.280 144.850 1303.540 145.170 ;
        RECT 1302.820 144.510 1303.080 144.830 ;
        RECT 1302.880 130.970 1303.020 144.510 ;
        RECT 1302.880 130.830 1303.480 130.970 ;
        RECT 1303.340 82.950 1303.480 130.830 ;
        RECT 1303.280 82.630 1303.540 82.950 ;
        RECT 1495.560 45.570 1495.820 45.890 ;
        RECT 1495.620 2.400 1495.760 45.570 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
      LAYER via2 ;
        RECT 1301.890 1621.320 1302.170 1621.600 ;
        RECT 1303.270 1621.320 1303.550 1621.600 ;
        RECT 1303.270 1332.320 1303.550 1332.600 ;
        RECT 1303.270 1331.640 1303.550 1331.920 ;
        RECT 1302.810 1138.520 1303.090 1138.800 ;
        RECT 1303.730 1138.520 1304.010 1138.800 ;
        RECT 1304.650 1041.960 1304.930 1042.240 ;
        RECT 1303.730 1041.280 1304.010 1041.560 ;
        RECT 1303.270 889.640 1303.550 889.920 ;
        RECT 1304.190 889.640 1304.470 889.920 ;
        RECT 1303.270 842.040 1303.550 842.320 ;
        RECT 1304.190 842.040 1304.470 842.320 ;
        RECT 1302.810 503.400 1303.090 503.680 ;
        RECT 1303.270 502.720 1303.550 503.000 ;
      LAYER met3 ;
        RECT 1301.865 1621.610 1302.195 1621.625 ;
        RECT 1303.245 1621.610 1303.575 1621.625 ;
        RECT 1301.865 1621.310 1303.575 1621.610 ;
        RECT 1301.865 1621.295 1302.195 1621.310 ;
        RECT 1303.245 1621.295 1303.575 1621.310 ;
        RECT 1303.245 1332.610 1303.575 1332.625 ;
        RECT 1303.030 1332.295 1303.575 1332.610 ;
        RECT 1303.030 1331.945 1303.330 1332.295 ;
        RECT 1303.030 1331.630 1303.575 1331.945 ;
        RECT 1303.245 1331.615 1303.575 1331.630 ;
        RECT 1302.785 1138.810 1303.115 1138.825 ;
        RECT 1303.705 1138.810 1304.035 1138.825 ;
        RECT 1302.785 1138.510 1304.035 1138.810 ;
        RECT 1302.785 1138.495 1303.115 1138.510 ;
        RECT 1303.705 1138.495 1304.035 1138.510 ;
        RECT 1304.625 1042.250 1304.955 1042.265 ;
        RECT 1303.950 1041.950 1304.955 1042.250 ;
        RECT 1303.950 1041.585 1304.250 1041.950 ;
        RECT 1304.625 1041.935 1304.955 1041.950 ;
        RECT 1303.705 1041.270 1304.250 1041.585 ;
        RECT 1303.705 1041.255 1304.035 1041.270 ;
        RECT 1303.245 889.930 1303.575 889.945 ;
        RECT 1304.165 889.930 1304.495 889.945 ;
        RECT 1303.245 889.630 1304.495 889.930 ;
        RECT 1303.245 889.615 1303.575 889.630 ;
        RECT 1304.165 889.615 1304.495 889.630 ;
        RECT 1303.245 842.330 1303.575 842.345 ;
        RECT 1304.165 842.330 1304.495 842.345 ;
        RECT 1303.245 842.030 1304.495 842.330 ;
        RECT 1303.245 842.015 1303.575 842.030 ;
        RECT 1304.165 842.015 1304.495 842.030 ;
        RECT 1302.785 503.690 1303.115 503.705 ;
        RECT 1302.785 503.375 1303.330 503.690 ;
        RECT 1303.030 503.025 1303.330 503.375 ;
        RECT 1303.030 502.710 1303.575 503.025 ;
        RECT 1303.245 502.695 1303.575 502.710 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1305.090 1683.920 1305.410 1683.980 ;
        RECT 1307.390 1683.920 1307.710 1683.980 ;
        RECT 1305.090 1683.780 1307.710 1683.920 ;
        RECT 1305.090 1683.720 1305.410 1683.780 ;
        RECT 1307.390 1683.720 1307.710 1683.780 ;
        RECT 1306.930 44.780 1307.250 44.840 ;
        RECT 1513.010 44.780 1513.330 44.840 ;
        RECT 1306.930 44.640 1513.330 44.780 ;
        RECT 1306.930 44.580 1307.250 44.640 ;
        RECT 1513.010 44.580 1513.330 44.640 ;
      LAYER via ;
        RECT 1305.120 1683.720 1305.380 1683.980 ;
        RECT 1307.420 1683.720 1307.680 1683.980 ;
        RECT 1306.960 44.580 1307.220 44.840 ;
        RECT 1513.040 44.580 1513.300 44.840 ;
      LAYER met2 ;
        RECT 1305.020 1700.340 1305.300 1704.000 ;
        RECT 1305.020 1700.000 1305.320 1700.340 ;
        RECT 1305.180 1684.010 1305.320 1700.000 ;
        RECT 1305.120 1683.690 1305.380 1684.010 ;
        RECT 1307.420 1683.690 1307.680 1684.010 ;
        RECT 1307.480 1632.410 1307.620 1683.690 ;
        RECT 1307.020 1632.270 1307.620 1632.410 ;
        RECT 1307.020 44.870 1307.160 1632.270 ;
        RECT 1306.960 44.550 1307.220 44.870 ;
        RECT 1513.040 44.550 1513.300 44.870 ;
        RECT 1513.100 2.400 1513.240 44.550 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 709.850 1625.440 710.170 1625.500 ;
        RECT 1223.670 1625.440 1223.990 1625.500 ;
        RECT 709.850 1625.300 1223.990 1625.440 ;
        RECT 709.850 1625.240 710.170 1625.300 ;
        RECT 1223.670 1625.240 1223.990 1625.300 ;
      LAYER via ;
        RECT 709.880 1625.240 710.140 1625.500 ;
        RECT 1223.700 1625.240 1223.960 1625.500 ;
      LAYER met2 ;
        RECT 1222.680 1700.340 1222.960 1704.000 ;
        RECT 1222.680 1700.000 1222.980 1700.340 ;
        RECT 1222.840 1664.370 1222.980 1700.000 ;
        RECT 1222.840 1664.230 1223.900 1664.370 ;
        RECT 1223.760 1625.530 1223.900 1664.230 ;
        RECT 709.880 1625.210 710.140 1625.530 ;
        RECT 1223.700 1625.210 1223.960 1625.530 ;
        RECT 709.940 24.210 710.080 1625.210 ;
        RECT 709.940 24.070 710.540 24.210 ;
        RECT 710.400 2.400 710.540 24.070 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1306.010 1664.880 1306.330 1664.940 ;
        RECT 1306.930 1664.880 1307.250 1664.940 ;
        RECT 1306.010 1664.740 1307.250 1664.880 ;
        RECT 1306.010 1664.680 1306.330 1664.740 ;
        RECT 1306.930 1664.680 1307.250 1664.740 ;
        RECT 1306.010 45.460 1306.330 45.520 ;
        RECT 1530.950 45.460 1531.270 45.520 ;
        RECT 1306.010 45.320 1531.270 45.460 ;
        RECT 1306.010 45.260 1306.330 45.320 ;
        RECT 1530.950 45.260 1531.270 45.320 ;
      LAYER via ;
        RECT 1306.040 1664.680 1306.300 1664.940 ;
        RECT 1306.960 1664.680 1307.220 1664.940 ;
        RECT 1306.040 45.260 1306.300 45.520 ;
        RECT 1530.980 45.260 1531.240 45.520 ;
      LAYER met2 ;
        RECT 1306.860 1700.340 1307.140 1704.000 ;
        RECT 1306.860 1700.000 1307.160 1700.340 ;
        RECT 1307.020 1664.970 1307.160 1700.000 ;
        RECT 1306.040 1664.650 1306.300 1664.970 ;
        RECT 1306.960 1664.650 1307.220 1664.970 ;
        RECT 1306.100 45.550 1306.240 1664.650 ;
        RECT 1306.040 45.230 1306.300 45.550 ;
        RECT 1530.980 45.230 1531.240 45.550 ;
        RECT 1531.040 2.400 1531.180 45.230 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1306.470 1666.580 1306.790 1666.640 ;
        RECT 1308.770 1666.580 1309.090 1666.640 ;
        RECT 1306.470 1666.440 1309.090 1666.580 ;
        RECT 1306.470 1666.380 1306.790 1666.440 ;
        RECT 1308.770 1666.380 1309.090 1666.440 ;
        RECT 1306.470 45.120 1306.790 45.180 ;
        RECT 1548.890 45.120 1549.210 45.180 ;
        RECT 1306.470 44.980 1549.210 45.120 ;
        RECT 1306.470 44.920 1306.790 44.980 ;
        RECT 1548.890 44.920 1549.210 44.980 ;
      LAYER via ;
        RECT 1306.500 1666.380 1306.760 1666.640 ;
        RECT 1308.800 1666.380 1309.060 1666.640 ;
        RECT 1306.500 44.920 1306.760 45.180 ;
        RECT 1548.920 44.920 1549.180 45.180 ;
      LAYER met2 ;
        RECT 1308.700 1700.340 1308.980 1704.000 ;
        RECT 1308.700 1700.000 1309.000 1700.340 ;
        RECT 1308.860 1666.670 1309.000 1700.000 ;
        RECT 1306.500 1666.350 1306.760 1666.670 ;
        RECT 1308.800 1666.350 1309.060 1666.670 ;
        RECT 1306.560 45.210 1306.700 1666.350 ;
        RECT 1306.500 44.890 1306.760 45.210 ;
        RECT 1548.920 44.890 1549.180 45.210 ;
        RECT 1548.980 2.400 1549.120 44.890 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1310.610 1654.340 1310.930 1654.400 ;
        RECT 1566.370 1654.340 1566.690 1654.400 ;
        RECT 1310.610 1654.200 1566.690 1654.340 ;
        RECT 1310.610 1654.140 1310.930 1654.200 ;
        RECT 1566.370 1654.140 1566.690 1654.200 ;
      LAYER via ;
        RECT 1310.640 1654.140 1310.900 1654.400 ;
        RECT 1566.400 1654.140 1566.660 1654.400 ;
      LAYER met2 ;
        RECT 1310.540 1700.340 1310.820 1704.000 ;
        RECT 1310.540 1700.000 1310.840 1700.340 ;
        RECT 1310.700 1654.430 1310.840 1700.000 ;
        RECT 1310.640 1654.110 1310.900 1654.430 ;
        RECT 1566.400 1654.110 1566.660 1654.430 ;
        RECT 1566.460 17.410 1566.600 1654.110 ;
        RECT 1566.460 17.270 1567.060 17.410 ;
        RECT 1566.920 2.400 1567.060 17.270 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1400.385 1668.125 1401.935 1668.295 ;
        RECT 1497.445 1668.125 1498.535 1668.295 ;
      LAYER mcon ;
        RECT 1401.765 1668.125 1401.935 1668.295 ;
        RECT 1498.365 1668.125 1498.535 1668.295 ;
      LAYER met1 ;
        RECT 1312.450 1685.960 1312.770 1686.020 ;
        RECT 1314.750 1685.960 1315.070 1686.020 ;
        RECT 1312.450 1685.820 1315.070 1685.960 ;
        RECT 1312.450 1685.760 1312.770 1685.820 ;
        RECT 1314.750 1685.760 1315.070 1685.820 ;
        RECT 1314.750 1668.280 1315.070 1668.340 ;
        RECT 1400.325 1668.280 1400.615 1668.325 ;
        RECT 1314.750 1668.140 1400.615 1668.280 ;
        RECT 1314.750 1668.080 1315.070 1668.140 ;
        RECT 1400.325 1668.095 1400.615 1668.140 ;
        RECT 1401.705 1668.280 1401.995 1668.325 ;
        RECT 1497.385 1668.280 1497.675 1668.325 ;
        RECT 1401.705 1668.140 1497.675 1668.280 ;
        RECT 1401.705 1668.095 1401.995 1668.140 ;
        RECT 1497.385 1668.095 1497.675 1668.140 ;
        RECT 1498.305 1668.280 1498.595 1668.325 ;
        RECT 1580.170 1668.280 1580.490 1668.340 ;
        RECT 1498.305 1668.140 1580.490 1668.280 ;
        RECT 1498.305 1668.095 1498.595 1668.140 ;
        RECT 1580.170 1668.080 1580.490 1668.140 ;
      LAYER via ;
        RECT 1312.480 1685.760 1312.740 1686.020 ;
        RECT 1314.780 1685.760 1315.040 1686.020 ;
        RECT 1314.780 1668.080 1315.040 1668.340 ;
        RECT 1580.200 1668.080 1580.460 1668.340 ;
      LAYER met2 ;
        RECT 1312.380 1700.340 1312.660 1704.000 ;
        RECT 1312.380 1700.000 1312.680 1700.340 ;
        RECT 1312.540 1686.050 1312.680 1700.000 ;
        RECT 1312.480 1685.730 1312.740 1686.050 ;
        RECT 1314.780 1685.730 1315.040 1686.050 ;
        RECT 1314.840 1668.370 1314.980 1685.730 ;
        RECT 1314.780 1668.050 1315.040 1668.370 ;
        RECT 1580.200 1668.050 1580.460 1668.370 ;
        RECT 1580.260 17.410 1580.400 1668.050 ;
        RECT 1580.260 17.270 1585.000 17.410 ;
        RECT 1584.860 2.400 1585.000 17.270 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1314.290 1684.260 1314.610 1684.320 ;
        RECT 1316.130 1684.260 1316.450 1684.320 ;
        RECT 1314.290 1684.120 1316.450 1684.260 ;
        RECT 1314.290 1684.060 1314.610 1684.120 ;
        RECT 1316.130 1684.060 1316.450 1684.120 ;
        RECT 1316.590 1633.600 1316.910 1633.660 ;
        RECT 1600.870 1633.600 1601.190 1633.660 ;
        RECT 1316.590 1633.460 1601.190 1633.600 ;
        RECT 1316.590 1633.400 1316.910 1633.460 ;
        RECT 1600.870 1633.400 1601.190 1633.460 ;
      LAYER via ;
        RECT 1314.320 1684.060 1314.580 1684.320 ;
        RECT 1316.160 1684.060 1316.420 1684.320 ;
        RECT 1316.620 1633.400 1316.880 1633.660 ;
        RECT 1600.900 1633.400 1601.160 1633.660 ;
      LAYER met2 ;
        RECT 1314.220 1700.340 1314.500 1704.000 ;
        RECT 1314.220 1700.000 1314.520 1700.340 ;
        RECT 1314.380 1684.350 1314.520 1700.000 ;
        RECT 1314.320 1684.030 1314.580 1684.350 ;
        RECT 1316.160 1684.030 1316.420 1684.350 ;
        RECT 1316.220 1656.890 1316.360 1684.030 ;
        RECT 1316.220 1656.750 1316.820 1656.890 ;
        RECT 1316.680 1633.690 1316.820 1656.750 ;
        RECT 1316.620 1633.370 1316.880 1633.690 ;
        RECT 1600.900 1633.370 1601.160 1633.690 ;
        RECT 1600.960 17.410 1601.100 1633.370 ;
        RECT 1600.960 17.270 1602.480 17.410 ;
        RECT 1602.340 2.400 1602.480 17.270 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1317.510 1647.200 1317.830 1647.260 ;
        RECT 1614.670 1647.200 1614.990 1647.260 ;
        RECT 1317.510 1647.060 1614.990 1647.200 ;
        RECT 1317.510 1647.000 1317.830 1647.060 ;
        RECT 1614.670 1647.000 1614.990 1647.060 ;
      LAYER via ;
        RECT 1317.540 1647.000 1317.800 1647.260 ;
        RECT 1614.700 1647.000 1614.960 1647.260 ;
      LAYER met2 ;
        RECT 1316.060 1700.410 1316.340 1704.000 ;
        RECT 1316.060 1700.270 1316.820 1700.410 ;
        RECT 1316.060 1700.000 1316.340 1700.270 ;
        RECT 1316.680 1678.140 1316.820 1700.270 ;
        RECT 1316.680 1678.000 1317.740 1678.140 ;
        RECT 1317.600 1647.290 1317.740 1678.000 ;
        RECT 1317.540 1646.970 1317.800 1647.290 ;
        RECT 1614.700 1646.970 1614.960 1647.290 ;
        RECT 1614.760 17.410 1614.900 1646.970 ;
        RECT 1614.760 17.270 1620.420 17.410 ;
        RECT 1620.280 2.400 1620.420 17.270 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1317.970 1692.080 1318.290 1692.140 ;
        RECT 1329.470 1692.080 1329.790 1692.140 ;
        RECT 1317.970 1691.940 1329.790 1692.080 ;
        RECT 1317.970 1691.880 1318.290 1691.940 ;
        RECT 1329.470 1691.880 1329.790 1691.940 ;
        RECT 1329.470 1674.740 1329.790 1674.800 ;
        RECT 1635.370 1674.740 1635.690 1674.800 ;
        RECT 1329.470 1674.600 1635.690 1674.740 ;
        RECT 1329.470 1674.540 1329.790 1674.600 ;
        RECT 1635.370 1674.540 1635.690 1674.600 ;
      LAYER via ;
        RECT 1318.000 1691.880 1318.260 1692.140 ;
        RECT 1329.500 1691.880 1329.760 1692.140 ;
        RECT 1329.500 1674.540 1329.760 1674.800 ;
        RECT 1635.400 1674.540 1635.660 1674.800 ;
      LAYER met2 ;
        RECT 1317.900 1700.340 1318.180 1704.000 ;
        RECT 1317.900 1700.000 1318.200 1700.340 ;
        RECT 1318.060 1692.170 1318.200 1700.000 ;
        RECT 1318.000 1691.850 1318.260 1692.170 ;
        RECT 1329.500 1691.850 1329.760 1692.170 ;
        RECT 1329.560 1674.830 1329.700 1691.850 ;
        RECT 1329.500 1674.510 1329.760 1674.830 ;
        RECT 1635.400 1674.510 1635.660 1674.830 ;
        RECT 1635.460 17.410 1635.600 1674.510 ;
        RECT 1635.460 17.270 1638.360 17.410 ;
        RECT 1638.220 2.400 1638.360 17.270 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1319.810 1689.700 1320.130 1689.760 ;
        RECT 1340.510 1689.700 1340.830 1689.760 ;
        RECT 1319.810 1689.560 1340.830 1689.700 ;
        RECT 1319.810 1689.500 1320.130 1689.560 ;
        RECT 1340.510 1689.500 1340.830 1689.560 ;
        RECT 1340.510 1681.880 1340.830 1681.940 ;
        RECT 1656.070 1681.880 1656.390 1681.940 ;
        RECT 1340.510 1681.740 1656.390 1681.880 ;
        RECT 1340.510 1681.680 1340.830 1681.740 ;
        RECT 1656.070 1681.680 1656.390 1681.740 ;
      LAYER via ;
        RECT 1319.840 1689.500 1320.100 1689.760 ;
        RECT 1340.540 1689.500 1340.800 1689.760 ;
        RECT 1340.540 1681.680 1340.800 1681.940 ;
        RECT 1656.100 1681.680 1656.360 1681.940 ;
      LAYER met2 ;
        RECT 1319.740 1700.340 1320.020 1704.000 ;
        RECT 1319.740 1700.000 1320.040 1700.340 ;
        RECT 1319.900 1689.790 1320.040 1700.000 ;
        RECT 1319.840 1689.470 1320.100 1689.790 ;
        RECT 1340.540 1689.470 1340.800 1689.790 ;
        RECT 1340.600 1681.970 1340.740 1689.470 ;
        RECT 1340.540 1681.650 1340.800 1681.970 ;
        RECT 1656.100 1681.650 1656.360 1681.970 ;
        RECT 1656.160 2.400 1656.300 1681.650 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1359.445 1660.985 1359.615 1662.175 ;
      LAYER mcon ;
        RECT 1359.445 1662.005 1359.615 1662.175 ;
      LAYER met1 ;
        RECT 1321.650 1686.640 1321.970 1686.700 ;
        RECT 1323.950 1686.640 1324.270 1686.700 ;
        RECT 1321.650 1686.500 1324.270 1686.640 ;
        RECT 1321.650 1686.440 1321.970 1686.500 ;
        RECT 1323.950 1686.440 1324.270 1686.500 ;
        RECT 1323.950 1662.160 1324.270 1662.220 ;
        RECT 1359.385 1662.160 1359.675 1662.205 ;
        RECT 1323.950 1662.020 1359.675 1662.160 ;
        RECT 1323.950 1661.960 1324.270 1662.020 ;
        RECT 1359.385 1661.975 1359.675 1662.020 ;
        RECT 1359.385 1661.140 1359.675 1661.185 ;
        RECT 1669.870 1661.140 1670.190 1661.200 ;
        RECT 1359.385 1661.000 1670.190 1661.140 ;
        RECT 1359.385 1660.955 1359.675 1661.000 ;
        RECT 1669.870 1660.940 1670.190 1661.000 ;
      LAYER via ;
        RECT 1321.680 1686.440 1321.940 1686.700 ;
        RECT 1323.980 1686.440 1324.240 1686.700 ;
        RECT 1323.980 1661.960 1324.240 1662.220 ;
        RECT 1669.900 1660.940 1670.160 1661.200 ;
      LAYER met2 ;
        RECT 1321.580 1700.340 1321.860 1704.000 ;
        RECT 1321.580 1700.000 1321.880 1700.340 ;
        RECT 1321.740 1686.730 1321.880 1700.000 ;
        RECT 1321.680 1686.410 1321.940 1686.730 ;
        RECT 1323.980 1686.410 1324.240 1686.730 ;
        RECT 1324.040 1662.250 1324.180 1686.410 ;
        RECT 1323.980 1661.930 1324.240 1662.250 ;
        RECT 1669.900 1660.910 1670.160 1661.230 ;
        RECT 1669.960 17.410 1670.100 1660.910 ;
        RECT 1669.960 17.270 1673.780 17.410 ;
        RECT 1673.640 2.400 1673.780 17.270 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1401.305 1667.785 1402.395 1667.955 ;
      LAYER mcon ;
        RECT 1402.225 1667.785 1402.395 1667.955 ;
      LAYER met1 ;
        RECT 1323.490 1667.940 1323.810 1668.000 ;
        RECT 1401.245 1667.940 1401.535 1667.985 ;
        RECT 1323.490 1667.800 1401.535 1667.940 ;
        RECT 1323.490 1667.740 1323.810 1667.800 ;
        RECT 1401.245 1667.755 1401.535 1667.800 ;
        RECT 1402.165 1667.940 1402.455 1667.985 ;
        RECT 1690.570 1667.940 1690.890 1668.000 ;
        RECT 1402.165 1667.800 1690.890 1667.940 ;
        RECT 1402.165 1667.755 1402.455 1667.800 ;
        RECT 1690.570 1667.740 1690.890 1667.800 ;
      LAYER via ;
        RECT 1323.520 1667.740 1323.780 1668.000 ;
        RECT 1690.600 1667.740 1690.860 1668.000 ;
      LAYER met2 ;
        RECT 1323.420 1700.340 1323.700 1704.000 ;
        RECT 1323.420 1700.000 1323.720 1700.340 ;
        RECT 1323.580 1668.030 1323.720 1700.000 ;
        RECT 1323.520 1667.710 1323.780 1668.030 ;
        RECT 1690.600 1667.710 1690.860 1668.030 ;
        RECT 1690.660 17.410 1690.800 1667.710 ;
        RECT 1690.660 17.270 1691.720 17.410 ;
        RECT 1691.580 2.400 1691.720 17.270 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1224.590 1678.140 1224.910 1678.200 ;
        RECT 1227.810 1678.140 1228.130 1678.200 ;
        RECT 1224.590 1678.000 1228.130 1678.140 ;
        RECT 1224.590 1677.940 1224.910 1678.000 ;
        RECT 1227.810 1677.940 1228.130 1678.000 ;
        RECT 731.010 1611.840 731.330 1611.900 ;
        RECT 1227.810 1611.840 1228.130 1611.900 ;
        RECT 731.010 1611.700 1228.130 1611.840 ;
        RECT 731.010 1611.640 731.330 1611.700 ;
        RECT 1227.810 1611.640 1228.130 1611.700 ;
      LAYER via ;
        RECT 1224.620 1677.940 1224.880 1678.200 ;
        RECT 1227.840 1677.940 1228.100 1678.200 ;
        RECT 731.040 1611.640 731.300 1611.900 ;
        RECT 1227.840 1611.640 1228.100 1611.900 ;
      LAYER met2 ;
        RECT 1224.520 1700.340 1224.800 1704.000 ;
        RECT 1224.520 1700.000 1224.820 1700.340 ;
        RECT 1224.680 1678.230 1224.820 1700.000 ;
        RECT 1224.620 1677.910 1224.880 1678.230 ;
        RECT 1227.840 1677.910 1228.100 1678.230 ;
        RECT 1227.900 1611.930 1228.040 1677.910 ;
        RECT 731.040 1611.610 731.300 1611.930 ;
        RECT 1227.840 1611.610 1228.100 1611.930 ;
        RECT 731.100 16.730 731.240 1611.610 ;
        RECT 728.340 16.590 731.240 16.730 ;
        RECT 728.340 2.400 728.480 16.590 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1325.330 50.220 1325.650 50.280 ;
        RECT 1704.370 50.220 1704.690 50.280 ;
        RECT 1325.330 50.080 1704.690 50.220 ;
        RECT 1325.330 50.020 1325.650 50.080 ;
        RECT 1704.370 50.020 1704.690 50.080 ;
      LAYER via ;
        RECT 1325.360 50.020 1325.620 50.280 ;
        RECT 1704.400 50.020 1704.660 50.280 ;
      LAYER met2 ;
        RECT 1325.260 1700.340 1325.540 1704.000 ;
        RECT 1325.260 1700.000 1325.560 1700.340 ;
        RECT 1325.420 50.310 1325.560 1700.000 ;
        RECT 1325.360 49.990 1325.620 50.310 ;
        RECT 1704.400 49.990 1704.660 50.310 ;
        RECT 1704.460 17.410 1704.600 49.990 ;
        RECT 1704.460 17.270 1709.660 17.410 ;
        RECT 1709.520 2.400 1709.660 17.270 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1327.170 1676.780 1327.490 1676.840 ;
        RECT 1327.630 1676.780 1327.950 1676.840 ;
        RECT 1327.170 1676.640 1327.950 1676.780 ;
        RECT 1327.170 1676.580 1327.490 1676.640 ;
        RECT 1327.630 1676.580 1327.950 1676.640 ;
        RECT 1327.630 1635.300 1327.950 1635.360 ;
        RECT 1328.090 1635.300 1328.410 1635.360 ;
        RECT 1327.630 1635.160 1328.410 1635.300 ;
        RECT 1327.630 1635.100 1327.950 1635.160 ;
        RECT 1328.090 1635.100 1328.410 1635.160 ;
        RECT 1328.550 50.560 1328.870 50.620 ;
        RECT 1725.070 50.560 1725.390 50.620 ;
        RECT 1328.550 50.420 1725.390 50.560 ;
        RECT 1328.550 50.360 1328.870 50.420 ;
        RECT 1725.070 50.360 1725.390 50.420 ;
      LAYER via ;
        RECT 1327.200 1676.580 1327.460 1676.840 ;
        RECT 1327.660 1676.580 1327.920 1676.840 ;
        RECT 1327.660 1635.100 1327.920 1635.360 ;
        RECT 1328.120 1635.100 1328.380 1635.360 ;
        RECT 1328.580 50.360 1328.840 50.620 ;
        RECT 1725.100 50.360 1725.360 50.620 ;
      LAYER met2 ;
        RECT 1327.100 1700.340 1327.380 1704.000 ;
        RECT 1327.100 1700.000 1327.400 1700.340 ;
        RECT 1327.260 1676.870 1327.400 1700.000 ;
        RECT 1327.200 1676.550 1327.460 1676.870 ;
        RECT 1327.660 1676.550 1327.920 1676.870 ;
        RECT 1327.720 1635.390 1327.860 1676.550 ;
        RECT 1327.660 1635.070 1327.920 1635.390 ;
        RECT 1328.120 1635.070 1328.380 1635.390 ;
        RECT 1328.180 1514.770 1328.320 1635.070 ;
        RECT 1328.180 1514.630 1328.780 1514.770 ;
        RECT 1328.640 50.650 1328.780 1514.630 ;
        RECT 1328.580 50.330 1328.840 50.650 ;
        RECT 1725.100 50.330 1725.360 50.650 ;
        RECT 1725.160 17.410 1725.300 50.330 ;
        RECT 1725.160 17.270 1727.600 17.410 ;
        RECT 1727.460 2.400 1727.600 17.270 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1329.010 50.900 1329.330 50.960 ;
        RECT 1738.870 50.900 1739.190 50.960 ;
        RECT 1329.010 50.760 1739.190 50.900 ;
        RECT 1329.010 50.700 1329.330 50.760 ;
        RECT 1738.870 50.700 1739.190 50.760 ;
        RECT 1738.870 20.980 1739.190 21.040 ;
        RECT 1745.310 20.980 1745.630 21.040 ;
        RECT 1738.870 20.840 1745.630 20.980 ;
        RECT 1738.870 20.780 1739.190 20.840 ;
        RECT 1745.310 20.780 1745.630 20.840 ;
      LAYER via ;
        RECT 1329.040 50.700 1329.300 50.960 ;
        RECT 1738.900 50.700 1739.160 50.960 ;
        RECT 1738.900 20.780 1739.160 21.040 ;
        RECT 1745.340 20.780 1745.600 21.040 ;
      LAYER met2 ;
        RECT 1328.940 1700.340 1329.220 1704.000 ;
        RECT 1328.940 1700.000 1329.240 1700.340 ;
        RECT 1329.100 50.990 1329.240 1700.000 ;
        RECT 1329.040 50.670 1329.300 50.990 ;
        RECT 1738.900 50.670 1739.160 50.990 ;
        RECT 1738.960 21.070 1739.100 50.670 ;
        RECT 1738.900 20.750 1739.160 21.070 ;
        RECT 1745.340 20.750 1745.600 21.070 ;
        RECT 1745.400 2.400 1745.540 20.750 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1329.930 51.240 1330.250 51.300 ;
        RECT 1759.570 51.240 1759.890 51.300 ;
        RECT 1329.930 51.100 1759.890 51.240 ;
        RECT 1329.930 51.040 1330.250 51.100 ;
        RECT 1759.570 51.040 1759.890 51.100 ;
      LAYER via ;
        RECT 1329.960 51.040 1330.220 51.300 ;
        RECT 1759.600 51.040 1759.860 51.300 ;
      LAYER met2 ;
        RECT 1330.780 1700.340 1331.060 1704.000 ;
        RECT 1330.780 1700.000 1331.080 1700.340 ;
        RECT 1330.940 1677.970 1331.080 1700.000 ;
        RECT 1330.020 1677.830 1331.080 1677.970 ;
        RECT 1330.020 51.330 1330.160 1677.830 ;
        RECT 1329.960 51.010 1330.220 51.330 ;
        RECT 1759.600 51.010 1759.860 51.330 ;
        RECT 1759.660 17.410 1759.800 51.010 ;
        RECT 1759.660 17.270 1763.020 17.410 ;
        RECT 1762.880 2.400 1763.020 17.270 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1337.365 1587.205 1337.535 1594.175 ;
        RECT 1337.365 331.245 1337.535 379.355 ;
      LAYER mcon ;
        RECT 1337.365 1594.005 1337.535 1594.175 ;
        RECT 1337.365 379.185 1337.535 379.355 ;
      LAYER met1 ;
        RECT 1332.690 1678.480 1333.010 1678.540 ;
        RECT 1337.290 1678.480 1337.610 1678.540 ;
        RECT 1332.690 1678.340 1337.610 1678.480 ;
        RECT 1332.690 1678.280 1333.010 1678.340 ;
        RECT 1337.290 1678.280 1337.610 1678.340 ;
        RECT 1337.290 1594.160 1337.610 1594.220 ;
        RECT 1337.095 1594.020 1337.610 1594.160 ;
        RECT 1337.290 1593.960 1337.610 1594.020 ;
        RECT 1337.290 1587.360 1337.610 1587.420 ;
        RECT 1337.095 1587.220 1337.610 1587.360 ;
        RECT 1337.290 1587.160 1337.610 1587.220 ;
        RECT 1337.290 379.340 1337.610 379.400 ;
        RECT 1337.095 379.200 1337.610 379.340 ;
        RECT 1337.290 379.140 1337.610 379.200 ;
        RECT 1337.290 331.400 1337.610 331.460 ;
        RECT 1337.095 331.260 1337.610 331.400 ;
        RECT 1337.290 331.200 1337.610 331.260 ;
        RECT 1337.290 54.980 1337.610 55.040 ;
        RECT 1780.730 54.980 1781.050 55.040 ;
        RECT 1337.290 54.840 1781.050 54.980 ;
        RECT 1337.290 54.780 1337.610 54.840 ;
        RECT 1780.730 54.780 1781.050 54.840 ;
      LAYER via ;
        RECT 1332.720 1678.280 1332.980 1678.540 ;
        RECT 1337.320 1678.280 1337.580 1678.540 ;
        RECT 1337.320 1593.960 1337.580 1594.220 ;
        RECT 1337.320 1587.160 1337.580 1587.420 ;
        RECT 1337.320 379.140 1337.580 379.400 ;
        RECT 1337.320 331.200 1337.580 331.460 ;
        RECT 1337.320 54.780 1337.580 55.040 ;
        RECT 1780.760 54.780 1781.020 55.040 ;
      LAYER met2 ;
        RECT 1332.620 1700.340 1332.900 1704.000 ;
        RECT 1332.620 1700.000 1332.920 1700.340 ;
        RECT 1332.780 1678.570 1332.920 1700.000 ;
        RECT 1332.720 1678.250 1332.980 1678.570 ;
        RECT 1337.320 1678.250 1337.580 1678.570 ;
        RECT 1337.380 1594.250 1337.520 1678.250 ;
        RECT 1337.320 1593.930 1337.580 1594.250 ;
        RECT 1337.320 1587.130 1337.580 1587.450 ;
        RECT 1337.380 379.430 1337.520 1587.130 ;
        RECT 1337.320 379.110 1337.580 379.430 ;
        RECT 1337.320 331.170 1337.580 331.490 ;
        RECT 1337.380 55.070 1337.520 331.170 ;
        RECT 1337.320 54.750 1337.580 55.070 ;
        RECT 1780.760 54.750 1781.020 55.070 ;
        RECT 1780.820 2.400 1780.960 54.750 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1334.530 1683.920 1334.850 1683.980 ;
        RECT 1336.830 1683.920 1337.150 1683.980 ;
        RECT 1334.530 1683.780 1337.150 1683.920 ;
        RECT 1334.530 1683.720 1334.850 1683.780 ;
        RECT 1336.830 1683.720 1337.150 1683.780 ;
        RECT 1336.370 54.640 1336.690 54.700 ;
        RECT 1794.070 54.640 1794.390 54.700 ;
        RECT 1336.370 54.500 1794.390 54.640 ;
        RECT 1336.370 54.440 1336.690 54.500 ;
        RECT 1794.070 54.440 1794.390 54.500 ;
      LAYER via ;
        RECT 1334.560 1683.720 1334.820 1683.980 ;
        RECT 1336.860 1683.720 1337.120 1683.980 ;
        RECT 1336.400 54.440 1336.660 54.700 ;
        RECT 1794.100 54.440 1794.360 54.700 ;
      LAYER met2 ;
        RECT 1334.460 1700.340 1334.740 1704.000 ;
        RECT 1334.460 1700.000 1334.760 1700.340 ;
        RECT 1334.620 1684.010 1334.760 1700.000 ;
        RECT 1334.560 1683.690 1334.820 1684.010 ;
        RECT 1336.860 1683.690 1337.120 1684.010 ;
        RECT 1336.920 1659.610 1337.060 1683.690 ;
        RECT 1336.460 1659.470 1337.060 1659.610 ;
        RECT 1336.460 54.730 1336.600 1659.470 ;
        RECT 1336.400 54.410 1336.660 54.730 ;
        RECT 1794.100 54.410 1794.360 54.730 ;
        RECT 1794.160 17.410 1794.300 54.410 ;
        RECT 1794.160 17.270 1798.900 17.410 ;
        RECT 1798.760 2.400 1798.900 17.270 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1335.910 54.300 1336.230 54.360 ;
        RECT 1814.770 54.300 1815.090 54.360 ;
        RECT 1335.910 54.160 1815.090 54.300 ;
        RECT 1335.910 54.100 1336.230 54.160 ;
        RECT 1814.770 54.100 1815.090 54.160 ;
      LAYER via ;
        RECT 1335.940 54.100 1336.200 54.360 ;
        RECT 1814.800 54.100 1815.060 54.360 ;
      LAYER met2 ;
        RECT 1336.300 1700.340 1336.580 1704.000 ;
        RECT 1336.300 1700.000 1336.600 1700.340 ;
        RECT 1336.460 1677.970 1336.600 1700.000 ;
        RECT 1336.000 1677.830 1336.600 1677.970 ;
        RECT 1336.000 54.390 1336.140 1677.830 ;
        RECT 1335.940 54.070 1336.200 54.390 ;
        RECT 1814.800 54.070 1815.060 54.390 ;
        RECT 1814.860 17.410 1815.000 54.070 ;
        RECT 1814.860 17.270 1816.840 17.410 ;
        RECT 1816.700 2.400 1816.840 17.270 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1336.830 1631.900 1337.150 1631.960 ;
        RECT 1338.210 1631.900 1338.530 1631.960 ;
        RECT 1336.830 1631.760 1338.530 1631.900 ;
        RECT 1336.830 1631.700 1337.150 1631.760 ;
        RECT 1338.210 1631.700 1338.530 1631.760 ;
        RECT 1336.830 53.960 1337.150 54.020 ;
        RECT 1828.570 53.960 1828.890 54.020 ;
        RECT 1336.830 53.820 1828.890 53.960 ;
        RECT 1336.830 53.760 1337.150 53.820 ;
        RECT 1828.570 53.760 1828.890 53.820 ;
        RECT 1828.570 20.980 1828.890 21.040 ;
        RECT 1834.550 20.980 1834.870 21.040 ;
        RECT 1828.570 20.840 1834.870 20.980 ;
        RECT 1828.570 20.780 1828.890 20.840 ;
        RECT 1834.550 20.780 1834.870 20.840 ;
      LAYER via ;
        RECT 1336.860 1631.700 1337.120 1631.960 ;
        RECT 1338.240 1631.700 1338.500 1631.960 ;
        RECT 1336.860 53.760 1337.120 54.020 ;
        RECT 1828.600 53.760 1828.860 54.020 ;
        RECT 1828.600 20.780 1828.860 21.040 ;
        RECT 1834.580 20.780 1834.840 21.040 ;
      LAYER met2 ;
        RECT 1338.140 1700.340 1338.420 1704.000 ;
        RECT 1338.140 1700.000 1338.440 1700.340 ;
        RECT 1338.300 1631.990 1338.440 1700.000 ;
        RECT 1336.860 1631.670 1337.120 1631.990 ;
        RECT 1338.240 1631.670 1338.500 1631.990 ;
        RECT 1336.920 54.050 1337.060 1631.670 ;
        RECT 1336.860 53.730 1337.120 54.050 ;
        RECT 1828.600 53.730 1828.860 54.050 ;
        RECT 1828.660 21.070 1828.800 53.730 ;
        RECT 1828.600 20.750 1828.860 21.070 ;
        RECT 1834.580 20.750 1834.840 21.070 ;
        RECT 1834.640 2.400 1834.780 20.750 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1345.185 1635.485 1345.355 1683.595 ;
        RECT 1344.265 841.925 1344.435 890.035 ;
        RECT 1344.265 752.165 1344.435 800.275 ;
        RECT 1344.265 559.385 1344.435 607.155 ;
        RECT 1344.265 503.625 1344.435 558.875 ;
        RECT 1344.265 435.285 1344.435 462.315 ;
        RECT 1344.725 358.785 1344.895 383.095 ;
        RECT 1344.265 83.045 1344.435 131.155 ;
      LAYER mcon ;
        RECT 1345.185 1683.425 1345.355 1683.595 ;
        RECT 1344.265 889.865 1344.435 890.035 ;
        RECT 1344.265 800.105 1344.435 800.275 ;
        RECT 1344.265 606.985 1344.435 607.155 ;
        RECT 1344.265 558.705 1344.435 558.875 ;
        RECT 1344.265 462.145 1344.435 462.315 ;
        RECT 1344.725 382.925 1344.895 383.095 ;
        RECT 1344.265 130.985 1344.435 131.155 ;
      LAYER met1 ;
        RECT 1340.050 1686.640 1340.370 1686.700 ;
        RECT 1345.110 1686.640 1345.430 1686.700 ;
        RECT 1340.050 1686.500 1345.430 1686.640 ;
        RECT 1340.050 1686.440 1340.370 1686.500 ;
        RECT 1345.110 1686.440 1345.430 1686.500 ;
        RECT 1345.110 1683.580 1345.430 1683.640 ;
        RECT 1344.915 1683.440 1345.430 1683.580 ;
        RECT 1345.110 1683.380 1345.430 1683.440 ;
        RECT 1345.110 1635.640 1345.430 1635.700 ;
        RECT 1344.915 1635.500 1345.430 1635.640 ;
        RECT 1345.110 1635.440 1345.430 1635.500 ;
        RECT 1344.190 1532.280 1344.510 1532.340 ;
        RECT 1345.110 1532.280 1345.430 1532.340 ;
        RECT 1344.190 1532.140 1345.430 1532.280 ;
        RECT 1344.190 1532.080 1344.510 1532.140 ;
        RECT 1345.110 1532.080 1345.430 1532.140 ;
        RECT 1344.190 1000.520 1344.510 1000.580 ;
        RECT 1345.110 1000.520 1345.430 1000.580 ;
        RECT 1344.190 1000.380 1345.430 1000.520 ;
        RECT 1344.190 1000.320 1344.510 1000.380 ;
        RECT 1345.110 1000.320 1345.430 1000.380 ;
        RECT 1344.190 890.020 1344.510 890.080 ;
        RECT 1343.995 889.880 1344.510 890.020 ;
        RECT 1344.190 889.820 1344.510 889.880 ;
        RECT 1344.205 842.080 1344.495 842.125 ;
        RECT 1344.650 842.080 1344.970 842.140 ;
        RECT 1344.205 841.940 1344.970 842.080 ;
        RECT 1344.205 841.895 1344.495 841.940 ;
        RECT 1344.650 841.880 1344.970 841.940 ;
        RECT 1344.190 807.400 1344.510 807.460 ;
        RECT 1344.650 807.400 1344.970 807.460 ;
        RECT 1344.190 807.260 1344.970 807.400 ;
        RECT 1344.190 807.200 1344.510 807.260 ;
        RECT 1344.650 807.200 1344.970 807.260 ;
        RECT 1344.190 800.260 1344.510 800.320 ;
        RECT 1343.995 800.120 1344.510 800.260 ;
        RECT 1344.190 800.060 1344.510 800.120 ;
        RECT 1344.205 752.320 1344.495 752.365 ;
        RECT 1344.650 752.320 1344.970 752.380 ;
        RECT 1344.205 752.180 1344.970 752.320 ;
        RECT 1344.205 752.135 1344.495 752.180 ;
        RECT 1344.650 752.120 1344.970 752.180 ;
        RECT 1344.190 710.840 1344.510 710.900 ;
        RECT 1344.650 710.840 1344.970 710.900 ;
        RECT 1344.190 710.700 1344.970 710.840 ;
        RECT 1344.190 710.640 1344.510 710.700 ;
        RECT 1344.650 710.640 1344.970 710.700 ;
        RECT 1344.190 607.140 1344.510 607.200 ;
        RECT 1343.995 607.000 1344.510 607.140 ;
        RECT 1344.190 606.940 1344.510 607.000 ;
        RECT 1344.190 559.540 1344.510 559.600 ;
        RECT 1343.995 559.400 1344.510 559.540 ;
        RECT 1344.190 559.340 1344.510 559.400 ;
        RECT 1344.190 558.860 1344.510 558.920 ;
        RECT 1343.995 558.720 1344.510 558.860 ;
        RECT 1344.190 558.660 1344.510 558.720 ;
        RECT 1344.190 503.780 1344.510 503.840 ;
        RECT 1343.995 503.640 1344.510 503.780 ;
        RECT 1344.190 503.580 1344.510 503.640 ;
        RECT 1344.190 462.300 1344.510 462.360 ;
        RECT 1343.995 462.160 1344.510 462.300 ;
        RECT 1344.190 462.100 1344.510 462.160 ;
        RECT 1344.205 435.440 1344.495 435.485 ;
        RECT 1344.650 435.440 1344.970 435.500 ;
        RECT 1344.205 435.300 1344.970 435.440 ;
        RECT 1344.205 435.255 1344.495 435.300 ;
        RECT 1344.650 435.240 1344.970 435.300 ;
        RECT 1344.650 383.080 1344.970 383.140 ;
        RECT 1344.455 382.940 1344.970 383.080 ;
        RECT 1344.650 382.880 1344.970 382.940 ;
        RECT 1344.665 358.940 1344.955 358.985 ;
        RECT 1345.110 358.940 1345.430 359.000 ;
        RECT 1344.665 358.800 1345.430 358.940 ;
        RECT 1344.665 358.755 1344.955 358.800 ;
        RECT 1345.110 358.740 1345.430 358.800 ;
        RECT 1344.190 342.620 1344.510 342.680 ;
        RECT 1345.110 342.620 1345.430 342.680 ;
        RECT 1344.190 342.480 1345.430 342.620 ;
        RECT 1344.190 342.420 1344.510 342.480 ;
        RECT 1345.110 342.420 1345.430 342.480 ;
        RECT 1344.190 131.140 1344.510 131.200 ;
        RECT 1343.995 131.000 1344.510 131.140 ;
        RECT 1344.190 130.940 1344.510 131.000 ;
        RECT 1344.190 83.200 1344.510 83.260 ;
        RECT 1343.995 83.060 1344.510 83.200 ;
        RECT 1344.190 83.000 1344.510 83.060 ;
        RECT 1344.190 53.620 1344.510 53.680 ;
        RECT 1849.270 53.620 1849.590 53.680 ;
        RECT 1344.190 53.480 1849.590 53.620 ;
        RECT 1344.190 53.420 1344.510 53.480 ;
        RECT 1849.270 53.420 1849.590 53.480 ;
      LAYER via ;
        RECT 1340.080 1686.440 1340.340 1686.700 ;
        RECT 1345.140 1686.440 1345.400 1686.700 ;
        RECT 1345.140 1683.380 1345.400 1683.640 ;
        RECT 1345.140 1635.440 1345.400 1635.700 ;
        RECT 1344.220 1532.080 1344.480 1532.340 ;
        RECT 1345.140 1532.080 1345.400 1532.340 ;
        RECT 1344.220 1000.320 1344.480 1000.580 ;
        RECT 1345.140 1000.320 1345.400 1000.580 ;
        RECT 1344.220 889.820 1344.480 890.080 ;
        RECT 1344.680 841.880 1344.940 842.140 ;
        RECT 1344.220 807.200 1344.480 807.460 ;
        RECT 1344.680 807.200 1344.940 807.460 ;
        RECT 1344.220 800.060 1344.480 800.320 ;
        RECT 1344.680 752.120 1344.940 752.380 ;
        RECT 1344.220 710.640 1344.480 710.900 ;
        RECT 1344.680 710.640 1344.940 710.900 ;
        RECT 1344.220 606.940 1344.480 607.200 ;
        RECT 1344.220 559.340 1344.480 559.600 ;
        RECT 1344.220 558.660 1344.480 558.920 ;
        RECT 1344.220 503.580 1344.480 503.840 ;
        RECT 1344.220 462.100 1344.480 462.360 ;
        RECT 1344.680 435.240 1344.940 435.500 ;
        RECT 1344.680 382.880 1344.940 383.140 ;
        RECT 1345.140 358.740 1345.400 359.000 ;
        RECT 1344.220 342.420 1344.480 342.680 ;
        RECT 1345.140 342.420 1345.400 342.680 ;
        RECT 1344.220 130.940 1344.480 131.200 ;
        RECT 1344.220 83.000 1344.480 83.260 ;
        RECT 1344.220 53.420 1344.480 53.680 ;
        RECT 1849.300 53.420 1849.560 53.680 ;
      LAYER met2 ;
        RECT 1339.980 1700.340 1340.260 1704.000 ;
        RECT 1339.980 1700.000 1340.280 1700.340 ;
        RECT 1340.140 1686.730 1340.280 1700.000 ;
        RECT 1340.080 1686.410 1340.340 1686.730 ;
        RECT 1345.140 1686.410 1345.400 1686.730 ;
        RECT 1345.200 1683.670 1345.340 1686.410 ;
        RECT 1345.140 1683.350 1345.400 1683.670 ;
        RECT 1345.140 1635.410 1345.400 1635.730 ;
        RECT 1345.200 1532.370 1345.340 1635.410 ;
        RECT 1344.220 1532.050 1344.480 1532.370 ;
        RECT 1345.140 1532.050 1345.400 1532.370 ;
        RECT 1344.280 1000.610 1344.420 1532.050 ;
        RECT 1344.220 1000.290 1344.480 1000.610 ;
        RECT 1345.140 1000.290 1345.400 1000.610 ;
        RECT 1345.200 952.525 1345.340 1000.290 ;
        RECT 1344.210 952.155 1344.490 952.525 ;
        RECT 1345.130 952.155 1345.410 952.525 ;
        RECT 1344.280 890.110 1344.420 952.155 ;
        RECT 1344.220 889.790 1344.480 890.110 ;
        RECT 1344.680 841.850 1344.940 842.170 ;
        RECT 1344.740 807.490 1344.880 841.850 ;
        RECT 1344.220 807.170 1344.480 807.490 ;
        RECT 1344.680 807.170 1344.940 807.490 ;
        RECT 1344.280 800.350 1344.420 807.170 ;
        RECT 1344.220 800.030 1344.480 800.350 ;
        RECT 1344.680 752.090 1344.940 752.410 ;
        RECT 1344.740 710.930 1344.880 752.090 ;
        RECT 1344.220 710.610 1344.480 710.930 ;
        RECT 1344.680 710.610 1344.940 710.930 ;
        RECT 1344.280 607.230 1344.420 710.610 ;
        RECT 1344.220 606.910 1344.480 607.230 ;
        RECT 1344.220 559.310 1344.480 559.630 ;
        RECT 1344.280 558.950 1344.420 559.310 ;
        RECT 1344.220 558.630 1344.480 558.950 ;
        RECT 1344.220 503.550 1344.480 503.870 ;
        RECT 1344.280 462.390 1344.420 503.550 ;
        RECT 1344.220 462.070 1344.480 462.390 ;
        RECT 1344.680 435.210 1344.940 435.530 ;
        RECT 1344.740 383.170 1344.880 435.210 ;
        RECT 1344.680 382.850 1344.940 383.170 ;
        RECT 1345.140 358.710 1345.400 359.030 ;
        RECT 1345.200 342.710 1345.340 358.710 ;
        RECT 1344.220 342.390 1344.480 342.710 ;
        RECT 1345.140 342.390 1345.400 342.710 ;
        RECT 1344.280 131.230 1344.420 342.390 ;
        RECT 1344.220 130.910 1344.480 131.230 ;
        RECT 1344.220 82.970 1344.480 83.290 ;
        RECT 1344.280 53.710 1344.420 82.970 ;
        RECT 1344.220 53.390 1344.480 53.710 ;
        RECT 1849.300 53.390 1849.560 53.710 ;
        RECT 1849.360 17.410 1849.500 53.390 ;
        RECT 1849.360 17.270 1852.260 17.410 ;
        RECT 1852.120 2.400 1852.260 17.270 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
      LAYER via2 ;
        RECT 1344.210 952.200 1344.490 952.480 ;
        RECT 1345.130 952.200 1345.410 952.480 ;
      LAYER met3 ;
        RECT 1344.185 952.490 1344.515 952.505 ;
        RECT 1345.105 952.490 1345.435 952.505 ;
        RECT 1344.185 952.190 1345.435 952.490 ;
        RECT 1344.185 952.175 1344.515 952.190 ;
        RECT 1345.105 952.175 1345.435 952.190 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1343.270 53.280 1343.590 53.340 ;
        RECT 1870.430 53.280 1870.750 53.340 ;
        RECT 1343.270 53.140 1870.750 53.280 ;
        RECT 1343.270 53.080 1343.590 53.140 ;
        RECT 1870.430 53.080 1870.750 53.140 ;
      LAYER via ;
        RECT 1343.300 53.080 1343.560 53.340 ;
        RECT 1870.460 53.080 1870.720 53.340 ;
      LAYER met2 ;
        RECT 1341.820 1700.410 1342.100 1704.000 ;
        RECT 1341.820 1700.270 1342.580 1700.410 ;
        RECT 1341.820 1700.000 1342.100 1700.270 ;
        RECT 1342.440 1677.970 1342.580 1700.270 ;
        RECT 1342.440 1677.830 1343.500 1677.970 ;
        RECT 1343.360 53.370 1343.500 1677.830 ;
        RECT 1343.300 53.050 1343.560 53.370 ;
        RECT 1870.460 53.050 1870.720 53.370 ;
        RECT 1870.520 7.210 1870.660 53.050 ;
        RECT 1870.060 7.070 1870.660 7.210 ;
        RECT 1870.060 2.400 1870.200 7.070 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 751.710 1605.040 752.030 1605.100 ;
        RECT 1225.970 1605.040 1226.290 1605.100 ;
        RECT 751.710 1604.900 1226.290 1605.040 ;
        RECT 751.710 1604.840 752.030 1604.900 ;
        RECT 1225.970 1604.840 1226.290 1604.900 ;
      LAYER via ;
        RECT 751.740 1604.840 752.000 1605.100 ;
        RECT 1226.000 1604.840 1226.260 1605.100 ;
      LAYER met2 ;
        RECT 1226.360 1700.340 1226.640 1704.000 ;
        RECT 1226.360 1700.000 1226.660 1700.340 ;
        RECT 1226.520 1616.770 1226.660 1700.000 ;
        RECT 1226.060 1616.630 1226.660 1616.770 ;
        RECT 1226.060 1605.130 1226.200 1616.630 ;
        RECT 751.740 1604.810 752.000 1605.130 ;
        RECT 1226.000 1604.810 1226.260 1605.130 ;
        RECT 751.800 16.730 751.940 1604.810 ;
        RECT 746.280 16.590 751.940 16.730 ;
        RECT 746.280 2.400 746.420 16.590 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1343.730 52.940 1344.050 53.000 ;
        RECT 1883.770 52.940 1884.090 53.000 ;
        RECT 1343.730 52.800 1884.090 52.940 ;
        RECT 1343.730 52.740 1344.050 52.800 ;
        RECT 1883.770 52.740 1884.090 52.800 ;
      LAYER via ;
        RECT 1343.760 52.740 1344.020 53.000 ;
        RECT 1883.800 52.740 1884.060 53.000 ;
      LAYER met2 ;
        RECT 1343.660 1700.340 1343.940 1704.000 ;
        RECT 1343.660 1700.000 1343.960 1700.340 ;
        RECT 1343.820 53.030 1343.960 1700.000 ;
        RECT 1343.760 52.710 1344.020 53.030 ;
        RECT 1883.800 52.710 1884.060 53.030 ;
        RECT 1883.860 17.410 1884.000 52.710 ;
        RECT 1883.860 17.270 1888.140 17.410 ;
        RECT 1888.000 2.400 1888.140 17.270 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1346.030 52.600 1346.350 52.660 ;
        RECT 1904.470 52.600 1904.790 52.660 ;
        RECT 1346.030 52.460 1904.790 52.600 ;
        RECT 1346.030 52.400 1346.350 52.460 ;
        RECT 1904.470 52.400 1904.790 52.460 ;
      LAYER via ;
        RECT 1346.060 52.400 1346.320 52.660 ;
        RECT 1904.500 52.400 1904.760 52.660 ;
      LAYER met2 ;
        RECT 1345.500 1700.410 1345.780 1704.000 ;
        RECT 1345.500 1700.270 1346.260 1700.410 ;
        RECT 1345.500 1700.000 1345.780 1700.270 ;
        RECT 1346.120 52.690 1346.260 1700.270 ;
        RECT 1346.060 52.370 1346.320 52.690 ;
        RECT 1904.500 52.370 1904.760 52.690 ;
        RECT 1904.560 17.410 1904.700 52.370 ;
        RECT 1904.560 17.270 1906.080 17.410 ;
        RECT 1905.940 2.400 1906.080 17.270 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1347.410 1684.600 1347.730 1684.660 ;
        RECT 1350.170 1684.600 1350.490 1684.660 ;
        RECT 1347.410 1684.460 1350.490 1684.600 ;
        RECT 1347.410 1684.400 1347.730 1684.460 ;
        RECT 1350.170 1684.400 1350.490 1684.460 ;
        RECT 1350.170 52.260 1350.490 52.320 ;
        RECT 1918.270 52.260 1918.590 52.320 ;
        RECT 1350.170 52.120 1918.590 52.260 ;
        RECT 1350.170 52.060 1350.490 52.120 ;
        RECT 1918.270 52.060 1918.590 52.120 ;
      LAYER via ;
        RECT 1347.440 1684.400 1347.700 1684.660 ;
        RECT 1350.200 1684.400 1350.460 1684.660 ;
        RECT 1350.200 52.060 1350.460 52.320 ;
        RECT 1918.300 52.060 1918.560 52.320 ;
      LAYER met2 ;
        RECT 1347.340 1700.340 1347.620 1704.000 ;
        RECT 1347.340 1700.000 1347.640 1700.340 ;
        RECT 1347.500 1684.690 1347.640 1700.000 ;
        RECT 1347.440 1684.370 1347.700 1684.690 ;
        RECT 1350.200 1684.370 1350.460 1684.690 ;
        RECT 1350.260 52.350 1350.400 1684.370 ;
        RECT 1350.200 52.030 1350.460 52.350 ;
        RECT 1918.300 52.030 1918.560 52.350 ;
        RECT 1918.360 17.410 1918.500 52.030 ;
        RECT 1918.360 17.270 1923.560 17.410 ;
        RECT 1923.420 2.400 1923.560 17.270 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1345.570 1685.280 1345.890 1685.340 ;
        RECT 1349.250 1685.280 1349.570 1685.340 ;
        RECT 1345.570 1685.140 1349.570 1685.280 ;
        RECT 1345.570 1685.080 1345.890 1685.140 ;
        RECT 1349.250 1685.080 1349.570 1685.140 ;
        RECT 1345.570 51.920 1345.890 51.980 ;
        RECT 1938.970 51.920 1939.290 51.980 ;
        RECT 1345.570 51.780 1939.290 51.920 ;
        RECT 1345.570 51.720 1345.890 51.780 ;
        RECT 1938.970 51.720 1939.290 51.780 ;
      LAYER via ;
        RECT 1345.600 1685.080 1345.860 1685.340 ;
        RECT 1349.280 1685.080 1349.540 1685.340 ;
        RECT 1345.600 51.720 1345.860 51.980 ;
        RECT 1939.000 51.720 1939.260 51.980 ;
      LAYER met2 ;
        RECT 1349.180 1700.340 1349.460 1704.000 ;
        RECT 1349.180 1700.000 1349.480 1700.340 ;
        RECT 1349.340 1685.370 1349.480 1700.000 ;
        RECT 1345.600 1685.050 1345.860 1685.370 ;
        RECT 1349.280 1685.050 1349.540 1685.370 ;
        RECT 1345.660 52.010 1345.800 1685.050 ;
        RECT 1345.600 51.690 1345.860 52.010 ;
        RECT 1939.000 51.690 1939.260 52.010 ;
        RECT 1939.060 17.410 1939.200 51.690 ;
        RECT 1939.060 17.270 1941.500 17.410 ;
        RECT 1941.360 2.400 1941.500 17.270 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1351.090 51.580 1351.410 51.640 ;
        RECT 1952.770 51.580 1953.090 51.640 ;
        RECT 1351.090 51.440 1953.090 51.580 ;
        RECT 1351.090 51.380 1351.410 51.440 ;
        RECT 1952.770 51.380 1953.090 51.440 ;
        RECT 1952.770 14.180 1953.090 14.240 ;
        RECT 1959.210 14.180 1959.530 14.240 ;
        RECT 1952.770 14.040 1959.530 14.180 ;
        RECT 1952.770 13.980 1953.090 14.040 ;
        RECT 1959.210 13.980 1959.530 14.040 ;
      LAYER via ;
        RECT 1351.120 51.380 1351.380 51.640 ;
        RECT 1952.800 51.380 1953.060 51.640 ;
        RECT 1952.800 13.980 1953.060 14.240 ;
        RECT 1959.240 13.980 1959.500 14.240 ;
      LAYER met2 ;
        RECT 1351.020 1700.340 1351.300 1704.000 ;
        RECT 1351.020 1700.000 1351.320 1700.340 ;
        RECT 1351.180 51.670 1351.320 1700.000 ;
        RECT 1351.120 51.350 1351.380 51.670 ;
        RECT 1952.800 51.350 1953.060 51.670 ;
        RECT 1952.860 14.270 1953.000 51.350 ;
        RECT 1952.800 13.950 1953.060 14.270 ;
        RECT 1959.240 13.950 1959.500 14.270 ;
        RECT 1959.300 2.400 1959.440 13.950 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.930 1605.380 1353.250 1605.440 ;
        RECT 1973.470 1605.380 1973.790 1605.440 ;
        RECT 1352.930 1605.240 1973.790 1605.380 ;
        RECT 1352.930 1605.180 1353.250 1605.240 ;
        RECT 1973.470 1605.180 1973.790 1605.240 ;
      LAYER via ;
        RECT 1352.960 1605.180 1353.220 1605.440 ;
        RECT 1973.500 1605.180 1973.760 1605.440 ;
      LAYER met2 ;
        RECT 1352.860 1700.340 1353.140 1704.000 ;
        RECT 1352.860 1700.000 1353.160 1700.340 ;
        RECT 1353.020 1605.470 1353.160 1700.000 ;
        RECT 1352.960 1605.150 1353.220 1605.470 ;
        RECT 1973.500 1605.150 1973.760 1605.470 ;
        RECT 1973.560 17.410 1973.700 1605.150 ;
        RECT 1973.560 17.270 1977.380 17.410 ;
        RECT 1977.240 2.400 1977.380 17.270 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1353.850 1625.780 1354.170 1625.840 ;
        RECT 1994.170 1625.780 1994.490 1625.840 ;
        RECT 1353.850 1625.640 1994.490 1625.780 ;
        RECT 1353.850 1625.580 1354.170 1625.640 ;
        RECT 1994.170 1625.580 1994.490 1625.640 ;
      LAYER via ;
        RECT 1353.880 1625.580 1354.140 1625.840 ;
        RECT 1994.200 1625.580 1994.460 1625.840 ;
      LAYER met2 ;
        RECT 1354.700 1700.340 1354.980 1704.000 ;
        RECT 1354.700 1700.000 1355.000 1700.340 ;
        RECT 1354.860 1661.650 1355.000 1700.000 ;
        RECT 1353.940 1661.510 1355.000 1661.650 ;
        RECT 1353.940 1625.870 1354.080 1661.510 ;
        RECT 1353.880 1625.550 1354.140 1625.870 ;
        RECT 1994.200 1625.550 1994.460 1625.870 ;
        RECT 1994.260 17.410 1994.400 1625.550 ;
        RECT 1994.260 17.270 1995.320 17.410 ;
        RECT 1995.180 2.400 1995.320 17.270 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1354.310 1661.140 1354.630 1661.200 ;
        RECT 1356.610 1661.140 1356.930 1661.200 ;
        RECT 1354.310 1661.000 1356.930 1661.140 ;
        RECT 1354.310 1660.940 1354.630 1661.000 ;
        RECT 1356.610 1660.940 1356.930 1661.000 ;
        RECT 1354.310 1591.100 1354.630 1591.160 ;
        RECT 2007.970 1591.100 2008.290 1591.160 ;
        RECT 1354.310 1590.960 2008.290 1591.100 ;
        RECT 1354.310 1590.900 1354.630 1590.960 ;
        RECT 2007.970 1590.900 2008.290 1590.960 ;
      LAYER via ;
        RECT 1354.340 1660.940 1354.600 1661.200 ;
        RECT 1356.640 1660.940 1356.900 1661.200 ;
        RECT 1354.340 1590.900 1354.600 1591.160 ;
        RECT 2008.000 1590.900 2008.260 1591.160 ;
      LAYER met2 ;
        RECT 1356.540 1700.340 1356.820 1704.000 ;
        RECT 1356.540 1700.000 1356.840 1700.340 ;
        RECT 1356.700 1661.230 1356.840 1700.000 ;
        RECT 1354.340 1660.910 1354.600 1661.230 ;
        RECT 1356.640 1660.910 1356.900 1661.230 ;
        RECT 1354.400 1591.190 1354.540 1660.910 ;
        RECT 1354.340 1590.870 1354.600 1591.190 ;
        RECT 2008.000 1590.870 2008.260 1591.190 ;
        RECT 2008.060 17.410 2008.200 1590.870 ;
        RECT 2008.060 17.270 2012.800 17.410 ;
        RECT 2012.660 2.400 2012.800 17.270 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1354.770 1660.800 1355.090 1660.860 ;
        RECT 1358.450 1660.800 1358.770 1660.860 ;
        RECT 1354.770 1660.660 1358.770 1660.800 ;
        RECT 1354.770 1660.600 1355.090 1660.660 ;
        RECT 1358.450 1660.600 1358.770 1660.660 ;
        RECT 1354.770 1535.680 1355.090 1535.740 ;
        RECT 2028.670 1535.680 2028.990 1535.740 ;
        RECT 1354.770 1535.540 2028.990 1535.680 ;
        RECT 1354.770 1535.480 1355.090 1535.540 ;
        RECT 2028.670 1535.480 2028.990 1535.540 ;
      LAYER via ;
        RECT 1354.800 1660.600 1355.060 1660.860 ;
        RECT 1358.480 1660.600 1358.740 1660.860 ;
        RECT 1354.800 1535.480 1355.060 1535.740 ;
        RECT 2028.700 1535.480 2028.960 1535.740 ;
      LAYER met2 ;
        RECT 1358.380 1700.340 1358.660 1704.000 ;
        RECT 1358.380 1700.000 1358.680 1700.340 ;
        RECT 1358.540 1660.890 1358.680 1700.000 ;
        RECT 1354.800 1660.570 1355.060 1660.890 ;
        RECT 1358.480 1660.570 1358.740 1660.890 ;
        RECT 1354.860 1535.770 1355.000 1660.570 ;
        RECT 1354.800 1535.450 1355.060 1535.770 ;
        RECT 2028.700 1535.450 2028.960 1535.770 ;
        RECT 2028.760 17.410 2028.900 1535.450 ;
        RECT 2028.760 17.270 2030.740 17.410 ;
        RECT 2030.600 2.400 2030.740 17.270 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1360.290 1584.300 1360.610 1584.360 ;
        RECT 2042.930 1584.300 2043.250 1584.360 ;
        RECT 1360.290 1584.160 2043.250 1584.300 ;
        RECT 1360.290 1584.100 1360.610 1584.160 ;
        RECT 2042.930 1584.100 2043.250 1584.160 ;
      LAYER via ;
        RECT 1360.320 1584.100 1360.580 1584.360 ;
        RECT 2042.960 1584.100 2043.220 1584.360 ;
      LAYER met2 ;
        RECT 1360.220 1700.340 1360.500 1704.000 ;
        RECT 1360.220 1700.000 1360.520 1700.340 ;
        RECT 1360.380 1584.390 1360.520 1700.000 ;
        RECT 1360.320 1584.070 1360.580 1584.390 ;
        RECT 2042.960 1584.070 2043.220 1584.390 ;
        RECT 2043.020 17.410 2043.160 1584.070 ;
        RECT 2043.020 17.270 2048.680 17.410 ;
        RECT 2048.540 2.400 2048.680 17.270 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 765.510 1660.460 765.830 1660.520 ;
        RECT 1228.270 1660.460 1228.590 1660.520 ;
        RECT 765.510 1660.320 1228.590 1660.460 ;
        RECT 765.510 1660.260 765.830 1660.320 ;
        RECT 1228.270 1660.260 1228.590 1660.320 ;
      LAYER via ;
        RECT 765.540 1660.260 765.800 1660.520 ;
        RECT 1228.300 1660.260 1228.560 1660.520 ;
      LAYER met2 ;
        RECT 1228.200 1700.340 1228.480 1704.000 ;
        RECT 1228.200 1700.000 1228.500 1700.340 ;
        RECT 1228.360 1660.550 1228.500 1700.000 ;
        RECT 765.540 1660.230 765.800 1660.550 ;
        RECT 1228.300 1660.230 1228.560 1660.550 ;
        RECT 765.600 18.090 765.740 1660.230 ;
        RECT 763.760 17.950 765.740 18.090 ;
        RECT 763.760 2.400 763.900 17.950 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1362.130 1528.540 1362.450 1528.600 ;
        RECT 2063.170 1528.540 2063.490 1528.600 ;
        RECT 1362.130 1528.400 2063.490 1528.540 ;
        RECT 1362.130 1528.340 1362.450 1528.400 ;
        RECT 2063.170 1528.340 2063.490 1528.400 ;
      LAYER via ;
        RECT 1362.160 1528.340 1362.420 1528.600 ;
        RECT 2063.200 1528.340 2063.460 1528.600 ;
      LAYER met2 ;
        RECT 1362.060 1700.340 1362.340 1704.000 ;
        RECT 1362.060 1700.000 1362.360 1700.340 ;
        RECT 1362.220 1528.630 1362.360 1700.000 ;
        RECT 1362.160 1528.310 1362.420 1528.630 ;
        RECT 2063.200 1528.310 2063.460 1528.630 ;
        RECT 2063.260 17.410 2063.400 1528.310 ;
        RECT 2063.260 17.270 2066.620 17.410 ;
        RECT 2066.480 2.400 2066.620 17.270 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1363.970 1459.520 1364.290 1459.580 ;
        RECT 2084.330 1459.520 2084.650 1459.580 ;
        RECT 1363.970 1459.380 2084.650 1459.520 ;
        RECT 1363.970 1459.320 1364.290 1459.380 ;
        RECT 2084.330 1459.320 2084.650 1459.380 ;
      LAYER via ;
        RECT 1364.000 1459.320 1364.260 1459.580 ;
        RECT 2084.360 1459.320 2084.620 1459.580 ;
      LAYER met2 ;
        RECT 1363.900 1700.340 1364.180 1704.000 ;
        RECT 1363.900 1700.000 1364.200 1700.340 ;
        RECT 1364.060 1459.610 1364.200 1700.000 ;
        RECT 1364.000 1459.290 1364.260 1459.610 ;
        RECT 2084.360 1459.290 2084.620 1459.610 ;
        RECT 2084.420 2.400 2084.560 1459.290 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1365.885 1635.485 1366.055 1683.595 ;
      LAYER mcon ;
        RECT 1365.885 1683.425 1366.055 1683.595 ;
      LAYER met1 ;
        RECT 1365.810 1683.580 1366.130 1683.640 ;
        RECT 1365.615 1683.440 1366.130 1683.580 ;
        RECT 1365.810 1683.380 1366.130 1683.440 ;
        RECT 1365.810 1635.640 1366.130 1635.700 ;
        RECT 1365.615 1635.500 1366.130 1635.640 ;
        RECT 1365.810 1635.440 1366.130 1635.500 ;
        RECT 1365.810 1521.740 1366.130 1521.800 ;
        RECT 2097.670 1521.740 2097.990 1521.800 ;
        RECT 1365.810 1521.600 2097.990 1521.740 ;
        RECT 1365.810 1521.540 1366.130 1521.600 ;
        RECT 2097.670 1521.540 2097.990 1521.600 ;
      LAYER via ;
        RECT 1365.840 1683.380 1366.100 1683.640 ;
        RECT 1365.840 1635.440 1366.100 1635.700 ;
        RECT 1365.840 1521.540 1366.100 1521.800 ;
        RECT 2097.700 1521.540 2097.960 1521.800 ;
      LAYER met2 ;
        RECT 1365.740 1700.340 1366.020 1704.000 ;
        RECT 1365.740 1700.000 1366.040 1700.340 ;
        RECT 1365.900 1683.670 1366.040 1700.000 ;
        RECT 1365.840 1683.350 1366.100 1683.670 ;
        RECT 1365.840 1635.410 1366.100 1635.730 ;
        RECT 1365.900 1521.830 1366.040 1635.410 ;
        RECT 1365.840 1521.510 1366.100 1521.830 ;
        RECT 2097.700 1521.510 2097.960 1521.830 ;
        RECT 2097.760 17.410 2097.900 1521.510 ;
        RECT 2097.760 17.270 2102.040 17.410 ;
        RECT 2101.900 2.400 2102.040 17.270 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1367.650 1684.940 1367.970 1685.000 ;
        RECT 1370.410 1684.940 1370.730 1685.000 ;
        RECT 1367.650 1684.800 1370.730 1684.940 ;
        RECT 1367.650 1684.740 1367.970 1684.800 ;
        RECT 1370.410 1684.740 1370.730 1684.800 ;
        RECT 1370.410 1577.160 1370.730 1577.220 ;
        RECT 2118.370 1577.160 2118.690 1577.220 ;
        RECT 1370.410 1577.020 2118.690 1577.160 ;
        RECT 1370.410 1576.960 1370.730 1577.020 ;
        RECT 2118.370 1576.960 2118.690 1577.020 ;
      LAYER via ;
        RECT 1367.680 1684.740 1367.940 1685.000 ;
        RECT 1370.440 1684.740 1370.700 1685.000 ;
        RECT 1370.440 1576.960 1370.700 1577.220 ;
        RECT 2118.400 1576.960 2118.660 1577.220 ;
      LAYER met2 ;
        RECT 1367.580 1700.340 1367.860 1704.000 ;
        RECT 1367.580 1700.000 1367.880 1700.340 ;
        RECT 1367.740 1685.030 1367.880 1700.000 ;
        RECT 1367.680 1684.710 1367.940 1685.030 ;
        RECT 1370.440 1684.710 1370.700 1685.030 ;
        RECT 1370.500 1577.250 1370.640 1684.710 ;
        RECT 1370.440 1576.930 1370.700 1577.250 ;
        RECT 2118.400 1576.930 2118.660 1577.250 ;
        RECT 2118.460 17.410 2118.600 1576.930 ;
        RECT 2118.460 17.270 2119.980 17.410 ;
        RECT 2119.840 2.400 2119.980 17.270 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1367.190 1683.920 1367.510 1683.980 ;
        RECT 1369.490 1683.920 1369.810 1683.980 ;
        RECT 1367.190 1683.780 1369.810 1683.920 ;
        RECT 1367.190 1683.720 1367.510 1683.780 ;
        RECT 1369.490 1683.720 1369.810 1683.780 ;
        RECT 1367.190 1514.940 1367.510 1515.000 ;
        RECT 2132.170 1514.940 2132.490 1515.000 ;
        RECT 1367.190 1514.800 2132.490 1514.940 ;
        RECT 1367.190 1514.740 1367.510 1514.800 ;
        RECT 2132.170 1514.740 2132.490 1514.800 ;
      LAYER via ;
        RECT 1367.220 1683.720 1367.480 1683.980 ;
        RECT 1369.520 1683.720 1369.780 1683.980 ;
        RECT 1367.220 1514.740 1367.480 1515.000 ;
        RECT 2132.200 1514.740 2132.460 1515.000 ;
      LAYER met2 ;
        RECT 1369.420 1700.340 1369.700 1704.000 ;
        RECT 1369.420 1700.000 1369.720 1700.340 ;
        RECT 1369.580 1684.010 1369.720 1700.000 ;
        RECT 1367.220 1683.690 1367.480 1684.010 ;
        RECT 1369.520 1683.690 1369.780 1684.010 ;
        RECT 1367.280 1515.030 1367.420 1683.690 ;
        RECT 1367.220 1514.710 1367.480 1515.030 ;
        RECT 2132.200 1514.710 2132.460 1515.030 ;
        RECT 2132.260 17.410 2132.400 1514.710 ;
        RECT 2132.260 17.270 2137.920 17.410 ;
        RECT 2137.780 2.400 2137.920 17.270 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1370.870 1452.720 1371.190 1452.780 ;
        RECT 2152.870 1452.720 2153.190 1452.780 ;
        RECT 1370.870 1452.580 2153.190 1452.720 ;
        RECT 1370.870 1452.520 1371.190 1452.580 ;
        RECT 2152.870 1452.520 2153.190 1452.580 ;
      LAYER via ;
        RECT 1370.900 1452.520 1371.160 1452.780 ;
        RECT 2152.900 1452.520 2153.160 1452.780 ;
      LAYER met2 ;
        RECT 1371.260 1700.340 1371.540 1704.000 ;
        RECT 1371.260 1700.000 1371.560 1700.340 ;
        RECT 1371.420 1631.900 1371.560 1700.000 ;
        RECT 1370.960 1631.760 1371.560 1631.900 ;
        RECT 1370.960 1452.810 1371.100 1631.760 ;
        RECT 1370.900 1452.490 1371.160 1452.810 ;
        RECT 2152.900 1452.490 2153.160 1452.810 ;
        RECT 2152.960 17.410 2153.100 1452.490 ;
        RECT 2152.960 17.270 2155.860 17.410 ;
        RECT 2155.720 2.400 2155.860 17.270 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1399.465 1632.425 1399.635 1633.955 ;
        RECT 1449.145 1632.425 1450.235 1632.595 ;
        RECT 1546.205 1632.425 1546.835 1632.595 ;
      LAYER mcon ;
        RECT 1399.465 1633.785 1399.635 1633.955 ;
        RECT 1450.065 1632.425 1450.235 1632.595 ;
        RECT 1546.665 1632.425 1546.835 1632.595 ;
      LAYER met1 ;
        RECT 1373.630 1633.940 1373.950 1634.000 ;
        RECT 1399.405 1633.940 1399.695 1633.985 ;
        RECT 1373.630 1633.800 1399.695 1633.940 ;
        RECT 1373.630 1633.740 1373.950 1633.800 ;
        RECT 1399.405 1633.755 1399.695 1633.800 ;
        RECT 1399.405 1632.580 1399.695 1632.625 ;
        RECT 1449.085 1632.580 1449.375 1632.625 ;
        RECT 1399.405 1632.440 1449.375 1632.580 ;
        RECT 1399.405 1632.395 1399.695 1632.440 ;
        RECT 1449.085 1632.395 1449.375 1632.440 ;
        RECT 1450.005 1632.580 1450.295 1632.625 ;
        RECT 1546.145 1632.580 1546.435 1632.625 ;
        RECT 1450.005 1632.440 1546.435 1632.580 ;
        RECT 1450.005 1632.395 1450.295 1632.440 ;
        RECT 1546.145 1632.395 1546.435 1632.440 ;
        RECT 1546.605 1632.580 1546.895 1632.625 ;
        RECT 2166.670 1632.580 2166.990 1632.640 ;
        RECT 1546.605 1632.440 2166.990 1632.580 ;
        RECT 1546.605 1632.395 1546.895 1632.440 ;
        RECT 2166.670 1632.380 2166.990 1632.440 ;
        RECT 2166.670 16.900 2166.990 16.960 ;
        RECT 2173.110 16.900 2173.430 16.960 ;
        RECT 2166.670 16.760 2173.430 16.900 ;
        RECT 2166.670 16.700 2166.990 16.760 ;
        RECT 2173.110 16.700 2173.430 16.760 ;
      LAYER via ;
        RECT 1373.660 1633.740 1373.920 1634.000 ;
        RECT 2166.700 1632.380 2166.960 1632.640 ;
        RECT 2166.700 16.700 2166.960 16.960 ;
        RECT 2173.140 16.700 2173.400 16.960 ;
      LAYER met2 ;
        RECT 1373.100 1700.410 1373.380 1704.000 ;
        RECT 1373.100 1700.270 1373.860 1700.410 ;
        RECT 1373.100 1700.000 1373.380 1700.270 ;
        RECT 1373.720 1634.030 1373.860 1700.270 ;
        RECT 1373.660 1633.710 1373.920 1634.030 ;
        RECT 2166.700 1632.350 2166.960 1632.670 ;
        RECT 2166.760 16.990 2166.900 1632.350 ;
        RECT 2166.700 16.670 2166.960 16.990 ;
        RECT 2173.140 16.670 2173.400 16.990 ;
        RECT 2173.200 2.400 2173.340 16.670 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1375.010 1683.920 1375.330 1683.980 ;
        RECT 1375.930 1683.920 1376.250 1683.980 ;
        RECT 1375.010 1683.780 1376.250 1683.920 ;
        RECT 1375.010 1683.720 1375.330 1683.780 ;
        RECT 1375.930 1683.720 1376.250 1683.780 ;
        RECT 1375.930 1618.640 1376.250 1618.700 ;
        RECT 2187.370 1618.640 2187.690 1618.700 ;
        RECT 1375.930 1618.500 2187.690 1618.640 ;
        RECT 1375.930 1618.440 1376.250 1618.500 ;
        RECT 2187.370 1618.440 2187.690 1618.500 ;
      LAYER via ;
        RECT 1375.040 1683.720 1375.300 1683.980 ;
        RECT 1375.960 1683.720 1376.220 1683.980 ;
        RECT 1375.960 1618.440 1376.220 1618.700 ;
        RECT 2187.400 1618.440 2187.660 1618.700 ;
      LAYER met2 ;
        RECT 1374.940 1700.340 1375.220 1704.000 ;
        RECT 1374.940 1700.000 1375.240 1700.340 ;
        RECT 1375.100 1684.010 1375.240 1700.000 ;
        RECT 1375.040 1683.690 1375.300 1684.010 ;
        RECT 1375.960 1683.690 1376.220 1684.010 ;
        RECT 1376.020 1618.730 1376.160 1683.690 ;
        RECT 1375.960 1618.410 1376.220 1618.730 ;
        RECT 2187.400 1618.410 2187.660 1618.730 ;
        RECT 2187.460 17.410 2187.600 1618.410 ;
        RECT 2187.460 17.270 2191.280 17.410 ;
        RECT 2191.140 2.400 2191.280 17.270 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1376.850 1570.360 1377.170 1570.420 ;
        RECT 2208.070 1570.360 2208.390 1570.420 ;
        RECT 1376.850 1570.220 2208.390 1570.360 ;
        RECT 1376.850 1570.160 1377.170 1570.220 ;
        RECT 2208.070 1570.160 2208.390 1570.220 ;
      LAYER via ;
        RECT 1376.880 1570.160 1377.140 1570.420 ;
        RECT 2208.100 1570.160 2208.360 1570.420 ;
      LAYER met2 ;
        RECT 1376.780 1700.340 1377.060 1704.000 ;
        RECT 1376.780 1700.000 1377.080 1700.340 ;
        RECT 1376.940 1570.450 1377.080 1700.000 ;
        RECT 1376.880 1570.130 1377.140 1570.450 ;
        RECT 2208.100 1570.130 2208.360 1570.450 ;
        RECT 2208.160 17.410 2208.300 1570.130 ;
        RECT 2208.160 17.270 2209.220 17.410 ;
        RECT 2209.080 2.400 2209.220 17.270 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1377.770 1507.800 1378.090 1507.860 ;
        RECT 2221.870 1507.800 2222.190 1507.860 ;
        RECT 1377.770 1507.660 2222.190 1507.800 ;
        RECT 1377.770 1507.600 1378.090 1507.660 ;
        RECT 2221.870 1507.600 2222.190 1507.660 ;
      LAYER via ;
        RECT 1377.800 1507.600 1378.060 1507.860 ;
        RECT 2221.900 1507.600 2222.160 1507.860 ;
      LAYER met2 ;
        RECT 1378.620 1700.340 1378.900 1704.000 ;
        RECT 1378.620 1700.000 1378.920 1700.340 ;
        RECT 1378.780 1665.730 1378.920 1700.000 ;
        RECT 1377.860 1665.590 1378.920 1665.730 ;
        RECT 1377.860 1507.890 1378.000 1665.590 ;
        RECT 1377.800 1507.570 1378.060 1507.890 ;
        RECT 2221.900 1507.570 2222.160 1507.890 ;
        RECT 2221.960 17.410 2222.100 1507.570 ;
        RECT 2221.960 17.270 2227.160 17.410 ;
        RECT 2227.020 2.400 2227.160 17.270 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 786.210 1646.520 786.530 1646.580 ;
        RECT 1230.110 1646.520 1230.430 1646.580 ;
        RECT 786.210 1646.380 1230.430 1646.520 ;
        RECT 786.210 1646.320 786.530 1646.380 ;
        RECT 1230.110 1646.320 1230.430 1646.380 ;
      LAYER via ;
        RECT 786.240 1646.320 786.500 1646.580 ;
        RECT 1230.140 1646.320 1230.400 1646.580 ;
      LAYER met2 ;
        RECT 1230.040 1700.340 1230.320 1704.000 ;
        RECT 1230.040 1700.000 1230.340 1700.340 ;
        RECT 1230.200 1646.610 1230.340 1700.000 ;
        RECT 786.240 1646.290 786.500 1646.610 ;
        RECT 1230.140 1646.290 1230.400 1646.610 ;
        RECT 786.300 18.090 786.440 1646.290 ;
        RECT 781.700 17.950 786.440 18.090 ;
        RECT 781.700 2.400 781.840 17.950 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1380.530 1666.580 1380.850 1666.640 ;
        RECT 1382.830 1666.580 1383.150 1666.640 ;
        RECT 1380.530 1666.440 1383.150 1666.580 ;
        RECT 1380.530 1666.380 1380.850 1666.440 ;
        RECT 1382.830 1666.380 1383.150 1666.440 ;
        RECT 1382.830 1605.040 1383.150 1605.100 ;
        RECT 2242.570 1605.040 2242.890 1605.100 ;
        RECT 1382.830 1604.900 2242.890 1605.040 ;
        RECT 1382.830 1604.840 1383.150 1604.900 ;
        RECT 2242.570 1604.840 2242.890 1604.900 ;
      LAYER via ;
        RECT 1380.560 1666.380 1380.820 1666.640 ;
        RECT 1382.860 1666.380 1383.120 1666.640 ;
        RECT 1382.860 1604.840 1383.120 1605.100 ;
        RECT 2242.600 1604.840 2242.860 1605.100 ;
      LAYER met2 ;
        RECT 1380.460 1700.340 1380.740 1704.000 ;
        RECT 1380.460 1700.000 1380.760 1700.340 ;
        RECT 1380.620 1666.670 1380.760 1700.000 ;
        RECT 1380.560 1666.350 1380.820 1666.670 ;
        RECT 1382.860 1666.350 1383.120 1666.670 ;
        RECT 1382.920 1605.130 1383.060 1666.350 ;
        RECT 1382.860 1604.810 1383.120 1605.130 ;
        RECT 2242.600 1604.810 2242.860 1605.130 ;
        RECT 2242.660 17.410 2242.800 1604.810 ;
        RECT 2242.660 17.270 2245.100 17.410 ;
        RECT 2244.960 2.400 2245.100 17.270 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1382.370 1683.920 1382.690 1683.980 ;
        RECT 1384.210 1683.920 1384.530 1683.980 ;
        RECT 1382.370 1683.780 1384.530 1683.920 ;
        RECT 1382.370 1683.720 1382.690 1683.780 ;
        RECT 1384.210 1683.720 1384.530 1683.780 ;
        RECT 1384.210 1445.920 1384.530 1445.980 ;
        RECT 2256.830 1445.920 2257.150 1445.980 ;
        RECT 1384.210 1445.780 2257.150 1445.920 ;
        RECT 1384.210 1445.720 1384.530 1445.780 ;
        RECT 2256.830 1445.720 2257.150 1445.780 ;
      LAYER via ;
        RECT 1382.400 1683.720 1382.660 1683.980 ;
        RECT 1384.240 1683.720 1384.500 1683.980 ;
        RECT 1384.240 1445.720 1384.500 1445.980 ;
        RECT 2256.860 1445.720 2257.120 1445.980 ;
      LAYER met2 ;
        RECT 1382.300 1700.340 1382.580 1704.000 ;
        RECT 1382.300 1700.000 1382.600 1700.340 ;
        RECT 1382.460 1684.010 1382.600 1700.000 ;
        RECT 1382.400 1683.690 1382.660 1684.010 ;
        RECT 1384.240 1683.690 1384.500 1684.010 ;
        RECT 1384.300 1446.010 1384.440 1683.690 ;
        RECT 1384.240 1445.690 1384.500 1446.010 ;
        RECT 2256.860 1445.690 2257.120 1446.010 ;
        RECT 2256.920 17.410 2257.060 1445.690 ;
        RECT 2256.920 17.270 2262.580 17.410 ;
        RECT 2262.440 2.400 2262.580 17.270 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1380.070 1684.940 1380.390 1685.000 ;
        RECT 1384.210 1684.940 1384.530 1685.000 ;
        RECT 1380.070 1684.800 1384.530 1684.940 ;
        RECT 1380.070 1684.740 1380.390 1684.800 ;
        RECT 1384.210 1684.740 1384.530 1684.800 ;
        RECT 1380.070 1501.000 1380.390 1501.060 ;
        RECT 2277.070 1501.000 2277.390 1501.060 ;
        RECT 1380.070 1500.860 2277.390 1501.000 ;
        RECT 1380.070 1500.800 1380.390 1500.860 ;
        RECT 2277.070 1500.800 2277.390 1500.860 ;
      LAYER via ;
        RECT 1380.100 1684.740 1380.360 1685.000 ;
        RECT 1384.240 1684.740 1384.500 1685.000 ;
        RECT 1380.100 1500.800 1380.360 1501.060 ;
        RECT 2277.100 1500.800 2277.360 1501.060 ;
      LAYER met2 ;
        RECT 1384.140 1700.340 1384.420 1704.000 ;
        RECT 1384.140 1700.000 1384.440 1700.340 ;
        RECT 1384.300 1685.030 1384.440 1700.000 ;
        RECT 1380.100 1684.710 1380.360 1685.030 ;
        RECT 1384.240 1684.710 1384.500 1685.030 ;
        RECT 1380.160 1501.090 1380.300 1684.710 ;
        RECT 1380.100 1500.770 1380.360 1501.090 ;
        RECT 2277.100 1500.770 2277.360 1501.090 ;
        RECT 2277.160 17.410 2277.300 1500.770 ;
        RECT 2277.160 17.270 2280.520 17.410 ;
        RECT 2280.380 2.400 2280.520 17.270 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1384.670 1686.980 1384.990 1687.040 ;
        RECT 1386.050 1686.980 1386.370 1687.040 ;
        RECT 1384.670 1686.840 1386.370 1686.980 ;
        RECT 1384.670 1686.780 1384.990 1686.840 ;
        RECT 1386.050 1686.780 1386.370 1686.840 ;
        RECT 1384.670 1438.440 1384.990 1438.500 ;
        RECT 2298.230 1438.440 2298.550 1438.500 ;
        RECT 1384.670 1438.300 2298.550 1438.440 ;
        RECT 1384.670 1438.240 1384.990 1438.300 ;
        RECT 2298.230 1438.240 2298.550 1438.300 ;
      LAYER via ;
        RECT 1384.700 1686.780 1384.960 1687.040 ;
        RECT 1386.080 1686.780 1386.340 1687.040 ;
        RECT 1384.700 1438.240 1384.960 1438.500 ;
        RECT 2298.260 1438.240 2298.520 1438.500 ;
      LAYER met2 ;
        RECT 1385.980 1700.340 1386.260 1704.000 ;
        RECT 1385.980 1700.000 1386.280 1700.340 ;
        RECT 1386.140 1687.070 1386.280 1700.000 ;
        RECT 1384.700 1686.750 1384.960 1687.070 ;
        RECT 1386.080 1686.750 1386.340 1687.070 ;
        RECT 1384.760 1438.530 1384.900 1686.750 ;
        RECT 1384.700 1438.210 1384.960 1438.530 ;
        RECT 2298.260 1438.210 2298.520 1438.530 ;
        RECT 2298.320 2.400 2298.460 1438.210 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1387.890 1684.940 1388.210 1685.000 ;
        RECT 1392.950 1684.940 1393.270 1685.000 ;
        RECT 1387.890 1684.800 1393.270 1684.940 ;
        RECT 1387.890 1684.740 1388.210 1684.800 ;
        RECT 1392.950 1684.740 1393.270 1684.800 ;
        RECT 1392.950 1652.980 1393.270 1653.040 ;
        RECT 2311.570 1652.980 2311.890 1653.040 ;
        RECT 1392.950 1652.840 2311.890 1652.980 ;
        RECT 1392.950 1652.780 1393.270 1652.840 ;
        RECT 2311.570 1652.780 2311.890 1652.840 ;
      LAYER via ;
        RECT 1387.920 1684.740 1388.180 1685.000 ;
        RECT 1392.980 1684.740 1393.240 1685.000 ;
        RECT 1392.980 1652.780 1393.240 1653.040 ;
        RECT 2311.600 1652.780 2311.860 1653.040 ;
      LAYER met2 ;
        RECT 1387.820 1700.340 1388.100 1704.000 ;
        RECT 1387.820 1700.000 1388.120 1700.340 ;
        RECT 1387.980 1685.030 1388.120 1700.000 ;
        RECT 1387.920 1684.710 1388.180 1685.030 ;
        RECT 1392.980 1684.710 1393.240 1685.030 ;
        RECT 1393.040 1653.070 1393.180 1684.710 ;
        RECT 1392.980 1652.750 1393.240 1653.070 ;
        RECT 2311.600 1652.750 2311.860 1653.070 ;
        RECT 2311.660 17.410 2311.800 1652.750 ;
        RECT 2311.660 17.270 2316.400 17.410 ;
        RECT 2316.260 2.400 2316.400 17.270 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1389.730 1683.920 1390.050 1683.980 ;
        RECT 1392.030 1683.920 1392.350 1683.980 ;
        RECT 1389.730 1683.780 1392.350 1683.920 ;
        RECT 1389.730 1683.720 1390.050 1683.780 ;
        RECT 1392.030 1683.720 1392.350 1683.780 ;
        RECT 1392.030 1563.560 1392.350 1563.620 ;
        RECT 2332.270 1563.560 2332.590 1563.620 ;
        RECT 1392.030 1563.420 2332.590 1563.560 ;
        RECT 1392.030 1563.360 1392.350 1563.420 ;
        RECT 2332.270 1563.360 2332.590 1563.420 ;
      LAYER via ;
        RECT 1389.760 1683.720 1390.020 1683.980 ;
        RECT 1392.060 1683.720 1392.320 1683.980 ;
        RECT 1392.060 1563.360 1392.320 1563.620 ;
        RECT 2332.300 1563.360 2332.560 1563.620 ;
      LAYER met2 ;
        RECT 1389.660 1700.340 1389.940 1704.000 ;
        RECT 1389.660 1700.000 1389.960 1700.340 ;
        RECT 1389.820 1684.010 1389.960 1700.000 ;
        RECT 1389.760 1683.690 1390.020 1684.010 ;
        RECT 1392.060 1683.690 1392.320 1684.010 ;
        RECT 1392.120 1563.650 1392.260 1683.690 ;
        RECT 1392.060 1563.330 1392.320 1563.650 ;
        RECT 2332.300 1563.330 2332.560 1563.650 ;
        RECT 2332.360 17.410 2332.500 1563.330 ;
        RECT 2332.360 17.270 2334.340 17.410 ;
        RECT 2334.200 2.400 2334.340 17.270 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1387.430 1684.260 1387.750 1684.320 ;
        RECT 1391.570 1684.260 1391.890 1684.320 ;
        RECT 1387.430 1684.120 1391.890 1684.260 ;
        RECT 1387.430 1684.060 1387.750 1684.120 ;
        RECT 1391.570 1684.060 1391.890 1684.120 ;
        RECT 1387.430 1611.500 1387.750 1611.560 ;
        RECT 2346.070 1611.500 2346.390 1611.560 ;
        RECT 1387.430 1611.360 2346.390 1611.500 ;
        RECT 1387.430 1611.300 1387.750 1611.360 ;
        RECT 2346.070 1611.300 2346.390 1611.360 ;
      LAYER via ;
        RECT 1387.460 1684.060 1387.720 1684.320 ;
        RECT 1391.600 1684.060 1391.860 1684.320 ;
        RECT 1387.460 1611.300 1387.720 1611.560 ;
        RECT 2346.100 1611.300 2346.360 1611.560 ;
      LAYER met2 ;
        RECT 1391.500 1700.340 1391.780 1704.000 ;
        RECT 1391.500 1700.000 1391.800 1700.340 ;
        RECT 1391.660 1684.350 1391.800 1700.000 ;
        RECT 1387.460 1684.030 1387.720 1684.350 ;
        RECT 1391.600 1684.030 1391.860 1684.350 ;
        RECT 1387.520 1611.590 1387.660 1684.030 ;
        RECT 1387.460 1611.270 1387.720 1611.590 ;
        RECT 2346.100 1611.270 2346.360 1611.590 ;
        RECT 2346.160 17.410 2346.300 1611.270 ;
        RECT 2346.160 17.270 2351.820 17.410 ;
        RECT 2351.680 2.400 2351.820 17.270 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1389.270 1685.280 1389.590 1685.340 ;
        RECT 1393.410 1685.280 1393.730 1685.340 ;
        RECT 1389.270 1685.140 1393.730 1685.280 ;
        RECT 1389.270 1685.080 1389.590 1685.140 ;
        RECT 1393.410 1685.080 1393.730 1685.140 ;
        RECT 1387.890 1683.920 1388.210 1683.980 ;
        RECT 1389.270 1683.920 1389.590 1683.980 ;
        RECT 1387.890 1683.780 1389.590 1683.920 ;
        RECT 1387.890 1683.720 1388.210 1683.780 ;
        RECT 1389.270 1683.720 1389.590 1683.780 ;
        RECT 1387.890 1493.860 1388.210 1493.920 ;
        RECT 2366.770 1493.860 2367.090 1493.920 ;
        RECT 1387.890 1493.720 2367.090 1493.860 ;
        RECT 1387.890 1493.660 1388.210 1493.720 ;
        RECT 2366.770 1493.660 2367.090 1493.720 ;
      LAYER via ;
        RECT 1389.300 1685.080 1389.560 1685.340 ;
        RECT 1393.440 1685.080 1393.700 1685.340 ;
        RECT 1387.920 1683.720 1388.180 1683.980 ;
        RECT 1389.300 1683.720 1389.560 1683.980 ;
        RECT 1387.920 1493.660 1388.180 1493.920 ;
        RECT 2366.800 1493.660 2367.060 1493.920 ;
      LAYER met2 ;
        RECT 1393.340 1700.340 1393.620 1704.000 ;
        RECT 1393.340 1700.000 1393.640 1700.340 ;
        RECT 1393.500 1685.370 1393.640 1700.000 ;
        RECT 1389.300 1685.050 1389.560 1685.370 ;
        RECT 1393.440 1685.050 1393.700 1685.370 ;
        RECT 1389.360 1684.010 1389.500 1685.050 ;
        RECT 1387.920 1683.690 1388.180 1684.010 ;
        RECT 1389.300 1683.690 1389.560 1684.010 ;
        RECT 1387.980 1493.950 1388.120 1683.690 ;
        RECT 1387.920 1493.630 1388.180 1493.950 ;
        RECT 2366.800 1493.630 2367.060 1493.950 ;
        RECT 2366.860 16.730 2367.000 1493.630 ;
        RECT 2366.860 16.590 2369.760 16.730 ;
        RECT 2369.620 2.400 2369.760 16.590 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1395.250 1677.460 1395.570 1677.520 ;
        RECT 1398.010 1677.460 1398.330 1677.520 ;
        RECT 1395.250 1677.320 1398.330 1677.460 ;
        RECT 1395.250 1677.260 1395.570 1677.320 ;
        RECT 1398.010 1677.260 1398.330 1677.320 ;
        RECT 1398.010 1431.640 1398.330 1431.700 ;
        RECT 2387.470 1431.640 2387.790 1431.700 ;
        RECT 1398.010 1431.500 2387.790 1431.640 ;
        RECT 1398.010 1431.440 1398.330 1431.500 ;
        RECT 2387.470 1431.440 2387.790 1431.500 ;
      LAYER via ;
        RECT 1395.280 1677.260 1395.540 1677.520 ;
        RECT 1398.040 1677.260 1398.300 1677.520 ;
        RECT 1398.040 1431.440 1398.300 1431.700 ;
        RECT 2387.500 1431.440 2387.760 1431.700 ;
      LAYER met2 ;
        RECT 1395.180 1700.340 1395.460 1704.000 ;
        RECT 1395.180 1700.000 1395.480 1700.340 ;
        RECT 1395.340 1677.550 1395.480 1700.000 ;
        RECT 1395.280 1677.230 1395.540 1677.550 ;
        RECT 1398.040 1677.230 1398.300 1677.550 ;
        RECT 1398.100 1431.730 1398.240 1677.230 ;
        RECT 1398.040 1431.410 1398.300 1431.730 ;
        RECT 2387.500 1431.410 2387.760 1431.730 ;
        RECT 2387.560 2.400 2387.700 1431.410 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1398.470 1424.840 1398.790 1424.900 ;
        RECT 2401.270 1424.840 2401.590 1424.900 ;
        RECT 1398.470 1424.700 2401.590 1424.840 ;
        RECT 1398.470 1424.640 1398.790 1424.700 ;
        RECT 2401.270 1424.640 2401.590 1424.700 ;
      LAYER via ;
        RECT 1398.500 1424.640 1398.760 1424.900 ;
        RECT 2401.300 1424.640 2401.560 1424.900 ;
      LAYER met2 ;
        RECT 1397.020 1700.340 1397.300 1704.000 ;
        RECT 1397.020 1700.000 1397.320 1700.340 ;
        RECT 1397.180 1677.970 1397.320 1700.000 ;
        RECT 1397.180 1677.830 1398.700 1677.970 ;
        RECT 1398.560 1424.930 1398.700 1677.830 ;
        RECT 1398.500 1424.610 1398.760 1424.930 ;
        RECT 2401.300 1424.610 2401.560 1424.930 ;
        RECT 2401.360 17.410 2401.500 1424.610 ;
        RECT 2401.360 17.270 2405.640 17.410 ;
        RECT 2405.500 2.400 2405.640 17.270 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 799.550 1632.580 799.870 1632.640 ;
        RECT 1231.950 1632.580 1232.270 1632.640 ;
        RECT 799.550 1632.440 1232.270 1632.580 ;
        RECT 799.550 1632.380 799.870 1632.440 ;
        RECT 1231.950 1632.380 1232.270 1632.440 ;
      LAYER via ;
        RECT 799.580 1632.380 799.840 1632.640 ;
        RECT 1231.980 1632.380 1232.240 1632.640 ;
      LAYER met2 ;
        RECT 1231.880 1700.340 1232.160 1704.000 ;
        RECT 1231.880 1700.000 1232.180 1700.340 ;
        RECT 1232.040 1632.670 1232.180 1700.000 ;
        RECT 799.580 1632.350 799.840 1632.670 ;
        RECT 1231.980 1632.350 1232.240 1632.670 ;
        RECT 799.640 2.400 799.780 1632.350 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1214.470 1679.160 1214.790 1679.220 ;
        RECT 1215.850 1679.160 1216.170 1679.220 ;
        RECT 1214.470 1679.020 1216.170 1679.160 ;
        RECT 1214.470 1678.960 1214.790 1679.020 ;
        RECT 1215.850 1678.960 1216.170 1679.020 ;
        RECT 648.210 1666.920 648.530 1666.980 ;
        RECT 1214.470 1666.920 1214.790 1666.980 ;
        RECT 648.210 1666.780 1214.790 1666.920 ;
        RECT 648.210 1666.720 648.530 1666.780 ;
        RECT 1214.470 1666.720 1214.790 1666.780 ;
      LAYER via ;
        RECT 1214.500 1678.960 1214.760 1679.220 ;
        RECT 1215.880 1678.960 1216.140 1679.220 ;
        RECT 648.240 1666.720 648.500 1666.980 ;
        RECT 1214.500 1666.720 1214.760 1666.980 ;
      LAYER met2 ;
        RECT 1215.780 1700.340 1216.060 1704.000 ;
        RECT 1215.780 1700.000 1216.080 1700.340 ;
        RECT 1215.940 1679.250 1216.080 1700.000 ;
        RECT 1214.500 1678.930 1214.760 1679.250 ;
        RECT 1215.880 1678.930 1216.140 1679.250 ;
        RECT 1214.560 1667.010 1214.700 1678.930 ;
        RECT 648.240 1666.690 648.500 1667.010 ;
        RECT 1214.500 1666.690 1214.760 1667.010 ;
        RECT 648.300 17.410 648.440 1666.690 ;
        RECT 645.080 17.270 648.440 17.410 ;
        RECT 645.080 2.400 645.220 17.270 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1396.630 1583.620 1396.950 1583.680 ;
        RECT 1398.930 1583.620 1399.250 1583.680 ;
        RECT 1396.630 1583.480 1399.250 1583.620 ;
        RECT 1396.630 1583.420 1396.950 1583.480 ;
        RECT 1398.930 1583.420 1399.250 1583.480 ;
        RECT 1396.630 1535.340 1396.950 1535.400 ;
        RECT 1398.930 1535.340 1399.250 1535.400 ;
        RECT 1396.630 1535.200 1399.250 1535.340 ;
        RECT 1396.630 1535.140 1396.950 1535.200 ;
        RECT 1398.930 1535.140 1399.250 1535.200 ;
        RECT 1398.930 1418.040 1399.250 1418.100 ;
        RECT 2428.870 1418.040 2429.190 1418.100 ;
        RECT 1398.930 1417.900 2429.190 1418.040 ;
        RECT 1398.930 1417.840 1399.250 1417.900 ;
        RECT 2428.870 1417.840 2429.190 1417.900 ;
      LAYER via ;
        RECT 1396.660 1583.420 1396.920 1583.680 ;
        RECT 1398.960 1583.420 1399.220 1583.680 ;
        RECT 1396.660 1535.140 1396.920 1535.400 ;
        RECT 1398.960 1535.140 1399.220 1535.400 ;
        RECT 1398.960 1417.840 1399.220 1418.100 ;
        RECT 2428.900 1417.840 2429.160 1418.100 ;
      LAYER met2 ;
        RECT 1399.320 1700.340 1399.600 1704.000 ;
        RECT 1399.320 1700.000 1399.620 1700.340 ;
        RECT 1399.480 1631.900 1399.620 1700.000 ;
        RECT 1399.020 1631.760 1399.620 1631.900 ;
        RECT 1399.020 1583.710 1399.160 1631.760 ;
        RECT 1396.660 1583.390 1396.920 1583.710 ;
        RECT 1398.960 1583.390 1399.220 1583.710 ;
        RECT 1396.720 1535.430 1396.860 1583.390 ;
        RECT 1396.660 1535.110 1396.920 1535.430 ;
        RECT 1398.960 1535.110 1399.220 1535.430 ;
        RECT 1399.020 1418.130 1399.160 1535.110 ;
        RECT 1398.960 1417.810 1399.220 1418.130 ;
        RECT 2428.900 1417.810 2429.160 1418.130 ;
        RECT 2428.960 2.400 2429.100 1417.810 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.770 1410.900 1401.090 1410.960 ;
        RECT 2442.670 1410.900 2442.990 1410.960 ;
        RECT 1400.770 1410.760 2442.990 1410.900 ;
        RECT 1400.770 1410.700 1401.090 1410.760 ;
        RECT 2442.670 1410.700 2442.990 1410.760 ;
      LAYER via ;
        RECT 1400.800 1410.700 1401.060 1410.960 ;
        RECT 2442.700 1410.700 2442.960 1410.960 ;
      LAYER met2 ;
        RECT 1401.160 1700.340 1401.440 1704.000 ;
        RECT 1401.160 1700.000 1401.460 1700.340 ;
        RECT 1401.320 1677.970 1401.460 1700.000 ;
        RECT 1400.860 1677.830 1401.460 1677.970 ;
        RECT 1400.860 1410.990 1401.000 1677.830 ;
        RECT 1400.800 1410.670 1401.060 1410.990 ;
        RECT 2442.700 1410.670 2442.960 1410.990 ;
        RECT 2442.760 18.090 2442.900 1410.670 ;
        RECT 2442.760 17.950 2447.040 18.090 ;
        RECT 2446.900 2.400 2447.040 17.950 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1403.070 1684.260 1403.390 1684.320 ;
        RECT 1406.750 1684.260 1407.070 1684.320 ;
        RECT 1403.070 1684.120 1407.070 1684.260 ;
        RECT 1403.070 1684.060 1403.390 1684.120 ;
        RECT 1406.750 1684.060 1407.070 1684.120 ;
        RECT 1406.290 1404.100 1406.610 1404.160 ;
        RECT 2463.370 1404.100 2463.690 1404.160 ;
        RECT 1406.290 1403.960 2463.690 1404.100 ;
        RECT 1406.290 1403.900 1406.610 1403.960 ;
        RECT 2463.370 1403.900 2463.690 1403.960 ;
        RECT 2463.370 2.960 2463.690 3.020 ;
        RECT 2464.750 2.960 2465.070 3.020 ;
        RECT 2463.370 2.820 2465.070 2.960 ;
        RECT 2463.370 2.760 2463.690 2.820 ;
        RECT 2464.750 2.760 2465.070 2.820 ;
      LAYER via ;
        RECT 1403.100 1684.060 1403.360 1684.320 ;
        RECT 1406.780 1684.060 1407.040 1684.320 ;
        RECT 1406.320 1403.900 1406.580 1404.160 ;
        RECT 2463.400 1403.900 2463.660 1404.160 ;
        RECT 2463.400 2.760 2463.660 3.020 ;
        RECT 2464.780 2.760 2465.040 3.020 ;
      LAYER met2 ;
        RECT 1403.000 1700.340 1403.280 1704.000 ;
        RECT 1403.000 1700.000 1403.300 1700.340 ;
        RECT 1403.160 1684.350 1403.300 1700.000 ;
        RECT 1403.100 1684.030 1403.360 1684.350 ;
        RECT 1406.780 1684.030 1407.040 1684.350 ;
        RECT 1406.840 1631.900 1406.980 1684.030 ;
        RECT 1406.380 1631.760 1406.980 1631.900 ;
        RECT 1406.380 1404.190 1406.520 1631.760 ;
        RECT 1406.320 1403.870 1406.580 1404.190 ;
        RECT 2463.400 1403.870 2463.660 1404.190 ;
        RECT 2463.460 3.050 2463.600 1403.870 ;
        RECT 2463.400 2.730 2463.660 3.050 ;
        RECT 2464.780 2.730 2465.040 3.050 ;
        RECT 2464.840 2.400 2464.980 2.730 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1404.910 1683.920 1405.230 1683.980 ;
        RECT 1407.210 1683.920 1407.530 1683.980 ;
        RECT 1404.910 1683.780 1407.530 1683.920 ;
        RECT 1404.910 1683.720 1405.230 1683.780 ;
        RECT 1407.210 1683.720 1407.530 1683.780 ;
        RECT 1406.750 1397.300 1407.070 1397.360 ;
        RECT 2477.170 1397.300 2477.490 1397.360 ;
        RECT 1406.750 1397.160 2477.490 1397.300 ;
        RECT 1406.750 1397.100 1407.070 1397.160 ;
        RECT 2477.170 1397.100 2477.490 1397.160 ;
        RECT 2477.170 2.960 2477.490 3.020 ;
        RECT 2482.690 2.960 2483.010 3.020 ;
        RECT 2477.170 2.820 2483.010 2.960 ;
        RECT 2477.170 2.760 2477.490 2.820 ;
        RECT 2482.690 2.760 2483.010 2.820 ;
      LAYER via ;
        RECT 1404.940 1683.720 1405.200 1683.980 ;
        RECT 1407.240 1683.720 1407.500 1683.980 ;
        RECT 1406.780 1397.100 1407.040 1397.360 ;
        RECT 2477.200 1397.100 2477.460 1397.360 ;
        RECT 2477.200 2.760 2477.460 3.020 ;
        RECT 2482.720 2.760 2482.980 3.020 ;
      LAYER met2 ;
        RECT 1404.840 1700.340 1405.120 1704.000 ;
        RECT 1404.840 1700.000 1405.140 1700.340 ;
        RECT 1405.000 1684.010 1405.140 1700.000 ;
        RECT 1404.940 1683.690 1405.200 1684.010 ;
        RECT 1407.240 1683.690 1407.500 1684.010 ;
        RECT 1407.300 1631.050 1407.440 1683.690 ;
        RECT 1406.840 1630.910 1407.440 1631.050 ;
        RECT 1406.840 1397.390 1406.980 1630.910 ;
        RECT 1406.780 1397.070 1407.040 1397.390 ;
        RECT 2477.200 1397.070 2477.460 1397.390 ;
        RECT 2477.260 3.050 2477.400 1397.070 ;
        RECT 2477.200 2.730 2477.460 3.050 ;
        RECT 2482.720 2.730 2482.980 3.050 ;
        RECT 2482.780 2.400 2482.920 2.730 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1403.530 1684.940 1403.850 1685.000 ;
        RECT 1406.750 1684.940 1407.070 1685.000 ;
        RECT 1403.530 1684.800 1407.070 1684.940 ;
        RECT 1403.530 1684.740 1403.850 1684.800 ;
        RECT 1406.750 1684.740 1407.070 1684.800 ;
        RECT 1401.690 1678.480 1402.010 1678.540 ;
        RECT 1403.530 1678.480 1403.850 1678.540 ;
        RECT 1401.690 1678.340 1403.850 1678.480 ;
        RECT 1401.690 1678.280 1402.010 1678.340 ;
        RECT 1403.530 1678.280 1403.850 1678.340 ;
        RECT 1401.230 1630.540 1401.550 1630.600 ;
        RECT 1407.210 1630.540 1407.530 1630.600 ;
        RECT 1401.230 1630.400 1407.530 1630.540 ;
        RECT 1401.230 1630.340 1401.550 1630.400 ;
        RECT 1407.210 1630.340 1407.530 1630.400 ;
        RECT 1407.210 900.560 1407.530 900.620 ;
        RECT 2497.870 900.560 2498.190 900.620 ;
        RECT 1407.210 900.420 2498.190 900.560 ;
        RECT 1407.210 900.360 1407.530 900.420 ;
        RECT 2497.870 900.360 2498.190 900.420 ;
      LAYER via ;
        RECT 1403.560 1684.740 1403.820 1685.000 ;
        RECT 1406.780 1684.740 1407.040 1685.000 ;
        RECT 1401.720 1678.280 1401.980 1678.540 ;
        RECT 1403.560 1678.280 1403.820 1678.540 ;
        RECT 1401.260 1630.340 1401.520 1630.600 ;
        RECT 1407.240 1630.340 1407.500 1630.600 ;
        RECT 1407.240 900.360 1407.500 900.620 ;
        RECT 2497.900 900.360 2498.160 900.620 ;
      LAYER met2 ;
        RECT 1406.680 1700.340 1406.960 1704.000 ;
        RECT 1406.680 1700.000 1406.980 1700.340 ;
        RECT 1406.840 1685.030 1406.980 1700.000 ;
        RECT 1403.560 1684.710 1403.820 1685.030 ;
        RECT 1406.780 1684.710 1407.040 1685.030 ;
        RECT 1403.620 1678.570 1403.760 1684.710 ;
        RECT 1401.720 1678.250 1401.980 1678.570 ;
        RECT 1403.560 1678.250 1403.820 1678.570 ;
        RECT 1401.780 1677.290 1401.920 1678.250 ;
        RECT 1401.320 1677.150 1401.920 1677.290 ;
        RECT 1401.320 1630.630 1401.460 1677.150 ;
        RECT 1401.260 1630.310 1401.520 1630.630 ;
        RECT 1407.240 1630.310 1407.500 1630.630 ;
        RECT 1407.300 900.650 1407.440 1630.310 ;
        RECT 1407.240 900.330 1407.500 900.650 ;
        RECT 2497.900 900.330 2498.160 900.650 ;
        RECT 2497.960 17.410 2498.100 900.330 ;
        RECT 2497.960 17.270 2500.860 17.410 ;
        RECT 2500.720 2.400 2500.860 17.270 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1408.590 1656.520 1408.910 1656.780 ;
        RECT 1408.680 1655.700 1408.820 1656.520 ;
        RECT 1424.690 1655.700 1425.010 1655.760 ;
        RECT 1408.680 1655.560 1425.010 1655.700 ;
        RECT 1424.690 1655.500 1425.010 1655.560 ;
        RECT 1424.690 1390.160 1425.010 1390.220 ;
        RECT 2512.130 1390.160 2512.450 1390.220 ;
        RECT 1424.690 1390.020 2512.450 1390.160 ;
        RECT 1424.690 1389.960 1425.010 1390.020 ;
        RECT 2512.130 1389.960 2512.450 1390.020 ;
        RECT 2512.130 18.260 2512.450 18.320 ;
        RECT 2518.110 18.260 2518.430 18.320 ;
        RECT 2512.130 18.120 2518.430 18.260 ;
        RECT 2512.130 18.060 2512.450 18.120 ;
        RECT 2518.110 18.060 2518.430 18.120 ;
      LAYER via ;
        RECT 1408.620 1656.520 1408.880 1656.780 ;
        RECT 1424.720 1655.500 1424.980 1655.760 ;
        RECT 1424.720 1389.960 1424.980 1390.220 ;
        RECT 2512.160 1389.960 2512.420 1390.220 ;
        RECT 2512.160 18.060 2512.420 18.320 ;
        RECT 2518.140 18.060 2518.400 18.320 ;
      LAYER met2 ;
        RECT 1408.520 1700.340 1408.800 1704.000 ;
        RECT 1408.520 1700.000 1408.820 1700.340 ;
        RECT 1408.680 1656.810 1408.820 1700.000 ;
        RECT 1408.620 1656.490 1408.880 1656.810 ;
        RECT 1424.720 1655.470 1424.980 1655.790 ;
        RECT 1424.780 1390.250 1424.920 1655.470 ;
        RECT 1424.720 1389.930 1424.980 1390.250 ;
        RECT 2512.160 1389.930 2512.420 1390.250 ;
        RECT 2512.220 18.350 2512.360 1389.930 ;
        RECT 2512.160 18.030 2512.420 18.350 ;
        RECT 2518.140 18.030 2518.400 18.350 ;
        RECT 2518.200 2.400 2518.340 18.030 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1410.430 1684.940 1410.750 1685.000 ;
        RECT 1413.190 1684.940 1413.510 1685.000 ;
        RECT 1410.430 1684.800 1413.510 1684.940 ;
        RECT 1410.430 1684.740 1410.750 1684.800 ;
        RECT 1413.190 1684.740 1413.510 1684.800 ;
        RECT 1413.190 1459.180 1413.510 1459.240 ;
        RECT 2532.370 1459.180 2532.690 1459.240 ;
        RECT 1413.190 1459.040 2532.690 1459.180 ;
        RECT 1413.190 1458.980 1413.510 1459.040 ;
        RECT 2532.370 1458.980 2532.690 1459.040 ;
      LAYER via ;
        RECT 1410.460 1684.740 1410.720 1685.000 ;
        RECT 1413.220 1684.740 1413.480 1685.000 ;
        RECT 1413.220 1458.980 1413.480 1459.240 ;
        RECT 2532.400 1458.980 2532.660 1459.240 ;
      LAYER met2 ;
        RECT 1410.360 1700.340 1410.640 1704.000 ;
        RECT 1410.360 1700.000 1410.660 1700.340 ;
        RECT 1410.520 1685.030 1410.660 1700.000 ;
        RECT 1410.460 1684.710 1410.720 1685.030 ;
        RECT 1413.220 1684.710 1413.480 1685.030 ;
        RECT 1413.280 1459.270 1413.420 1684.710 ;
        RECT 1413.220 1458.950 1413.480 1459.270 ;
        RECT 2532.400 1458.950 2532.660 1459.270 ;
        RECT 2532.460 17.410 2532.600 1458.950 ;
        RECT 2532.460 17.270 2536.280 17.410 ;
        RECT 2536.140 2.400 2536.280 17.270 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1409.510 1684.260 1409.830 1684.320 ;
        RECT 1412.270 1684.260 1412.590 1684.320 ;
        RECT 1409.510 1684.120 1412.590 1684.260 ;
        RECT 1409.510 1684.060 1409.830 1684.120 ;
        RECT 1412.270 1684.060 1412.590 1684.120 ;
        RECT 1409.970 1383.360 1410.290 1383.420 ;
        RECT 2553.070 1383.360 2553.390 1383.420 ;
        RECT 1409.970 1383.220 2553.390 1383.360 ;
        RECT 1409.970 1383.160 1410.290 1383.220 ;
        RECT 2553.070 1383.160 2553.390 1383.220 ;
      LAYER via ;
        RECT 1409.540 1684.060 1409.800 1684.320 ;
        RECT 1412.300 1684.060 1412.560 1684.320 ;
        RECT 1410.000 1383.160 1410.260 1383.420 ;
        RECT 2553.100 1383.160 2553.360 1383.420 ;
      LAYER met2 ;
        RECT 1412.200 1700.340 1412.480 1704.000 ;
        RECT 1412.200 1700.000 1412.500 1700.340 ;
        RECT 1412.360 1684.350 1412.500 1700.000 ;
        RECT 1409.540 1684.030 1409.800 1684.350 ;
        RECT 1412.300 1684.030 1412.560 1684.350 ;
        RECT 1409.600 1667.770 1409.740 1684.030 ;
        RECT 1409.600 1667.630 1410.200 1667.770 ;
        RECT 1410.060 1383.450 1410.200 1667.630 ;
        RECT 1410.000 1383.130 1410.260 1383.450 ;
        RECT 2553.100 1383.130 2553.360 1383.450 ;
        RECT 2553.160 17.410 2553.300 1383.130 ;
        RECT 2553.160 17.270 2554.220 17.410 ;
        RECT 2554.080 2.400 2554.220 17.270 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1411.350 1684.600 1411.670 1684.660 ;
        RECT 1414.110 1684.600 1414.430 1684.660 ;
        RECT 1411.350 1684.460 1414.430 1684.600 ;
        RECT 1411.350 1684.400 1411.670 1684.460 ;
        RECT 1414.110 1684.400 1414.430 1684.460 ;
        RECT 1411.350 1369.760 1411.670 1369.820 ;
        RECT 2566.870 1369.760 2567.190 1369.820 ;
        RECT 1411.350 1369.620 2567.190 1369.760 ;
        RECT 1411.350 1369.560 1411.670 1369.620 ;
        RECT 2566.870 1369.560 2567.190 1369.620 ;
      LAYER via ;
        RECT 1411.380 1684.400 1411.640 1684.660 ;
        RECT 1414.140 1684.400 1414.400 1684.660 ;
        RECT 1411.380 1369.560 1411.640 1369.820 ;
        RECT 2566.900 1369.560 2567.160 1369.820 ;
      LAYER met2 ;
        RECT 1414.040 1700.340 1414.320 1704.000 ;
        RECT 1414.040 1700.000 1414.340 1700.340 ;
        RECT 1414.200 1684.690 1414.340 1700.000 ;
        RECT 1411.380 1684.370 1411.640 1684.690 ;
        RECT 1414.140 1684.370 1414.400 1684.690 ;
        RECT 1411.440 1369.850 1411.580 1684.370 ;
        RECT 1411.380 1369.530 1411.640 1369.850 ;
        RECT 2566.900 1369.530 2567.160 1369.850 ;
        RECT 2566.960 17.410 2567.100 1369.530 ;
        RECT 2566.960 17.270 2572.160 17.410 ;
        RECT 2572.020 2.400 2572.160 17.270 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1415.030 1362.620 1415.350 1362.680 ;
        RECT 2587.570 1362.620 2587.890 1362.680 ;
        RECT 1415.030 1362.480 2587.890 1362.620 ;
        RECT 1415.030 1362.420 1415.350 1362.480 ;
        RECT 2587.570 1362.420 2587.890 1362.480 ;
      LAYER via ;
        RECT 1415.060 1362.420 1415.320 1362.680 ;
        RECT 2587.600 1362.420 2587.860 1362.680 ;
      LAYER met2 ;
        RECT 1415.880 1700.340 1416.160 1704.000 ;
        RECT 1415.880 1700.000 1416.180 1700.340 ;
        RECT 1416.040 1677.970 1416.180 1700.000 ;
        RECT 1415.120 1677.830 1416.180 1677.970 ;
        RECT 1415.120 1362.710 1415.260 1677.830 ;
        RECT 1415.060 1362.390 1415.320 1362.710 ;
        RECT 2587.600 1362.390 2587.860 1362.710 ;
        RECT 2587.660 17.410 2587.800 1362.390 ;
        RECT 2587.660 17.270 2589.640 17.410 ;
        RECT 2589.500 2.400 2589.640 17.270 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1229.650 1678.140 1229.970 1678.200 ;
        RECT 1234.250 1678.140 1234.570 1678.200 ;
        RECT 1229.650 1678.000 1234.570 1678.140 ;
        RECT 1229.650 1677.940 1229.970 1678.000 ;
        RECT 1234.250 1677.940 1234.570 1678.000 ;
        RECT 827.610 1618.640 827.930 1618.700 ;
        RECT 1229.650 1618.640 1229.970 1618.700 ;
        RECT 827.610 1618.500 1229.970 1618.640 ;
        RECT 827.610 1618.440 827.930 1618.500 ;
        RECT 1229.650 1618.440 1229.970 1618.500 ;
      LAYER via ;
        RECT 1229.680 1677.940 1229.940 1678.200 ;
        RECT 1234.280 1677.940 1234.540 1678.200 ;
        RECT 827.640 1618.440 827.900 1618.700 ;
        RECT 1229.680 1618.440 1229.940 1618.700 ;
      LAYER met2 ;
        RECT 1234.180 1700.340 1234.460 1704.000 ;
        RECT 1234.180 1700.000 1234.480 1700.340 ;
        RECT 1234.340 1678.230 1234.480 1700.000 ;
        RECT 1229.680 1677.910 1229.940 1678.230 ;
        RECT 1234.280 1677.910 1234.540 1678.230 ;
        RECT 1229.740 1618.730 1229.880 1677.910 ;
        RECT 827.640 1618.410 827.900 1618.730 ;
        RECT 1229.680 1618.410 1229.940 1618.730 ;
        RECT 827.700 17.410 827.840 1618.410 ;
        RECT 823.560 17.270 827.840 17.410 ;
        RECT 823.560 2.400 823.700 17.270 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1417.790 1677.120 1418.110 1677.180 ;
        RECT 1420.550 1677.120 1420.870 1677.180 ;
        RECT 1417.790 1676.980 1420.870 1677.120 ;
        RECT 1417.790 1676.920 1418.110 1676.980 ;
        RECT 1420.550 1676.920 1420.870 1676.980 ;
        RECT 1420.550 1355.820 1420.870 1355.880 ;
        RECT 2601.830 1355.820 2602.150 1355.880 ;
        RECT 1420.550 1355.680 2602.150 1355.820 ;
        RECT 1420.550 1355.620 1420.870 1355.680 ;
        RECT 2601.830 1355.620 2602.150 1355.680 ;
      LAYER via ;
        RECT 1417.820 1676.920 1418.080 1677.180 ;
        RECT 1420.580 1676.920 1420.840 1677.180 ;
        RECT 1420.580 1355.620 1420.840 1355.880 ;
        RECT 2601.860 1355.620 2602.120 1355.880 ;
      LAYER met2 ;
        RECT 1417.720 1700.340 1418.000 1704.000 ;
        RECT 1417.720 1700.000 1418.020 1700.340 ;
        RECT 1417.880 1677.210 1418.020 1700.000 ;
        RECT 1417.820 1676.890 1418.080 1677.210 ;
        RECT 1420.580 1676.890 1420.840 1677.210 ;
        RECT 1420.640 1355.910 1420.780 1676.890 ;
        RECT 1420.580 1355.590 1420.840 1355.910 ;
        RECT 2601.860 1355.590 2602.120 1355.910 ;
        RECT 2601.920 17.410 2602.060 1355.590 ;
        RECT 2601.920 17.270 2607.580 17.410 ;
        RECT 2607.440 2.400 2607.580 17.270 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1416.410 1684.260 1416.730 1684.320 ;
        RECT 1419.630 1684.260 1419.950 1684.320 ;
        RECT 1416.410 1684.120 1419.950 1684.260 ;
        RECT 1416.410 1684.060 1416.730 1684.120 ;
        RECT 1419.630 1684.060 1419.950 1684.120 ;
        RECT 1415.950 1349.020 1416.270 1349.080 ;
        RECT 2622.070 1349.020 2622.390 1349.080 ;
        RECT 1415.950 1348.880 2622.390 1349.020 ;
        RECT 1415.950 1348.820 1416.270 1348.880 ;
        RECT 2622.070 1348.820 2622.390 1348.880 ;
      LAYER via ;
        RECT 1416.440 1684.060 1416.700 1684.320 ;
        RECT 1419.660 1684.060 1419.920 1684.320 ;
        RECT 1415.980 1348.820 1416.240 1349.080 ;
        RECT 2622.100 1348.820 2622.360 1349.080 ;
      LAYER met2 ;
        RECT 1419.560 1700.340 1419.840 1704.000 ;
        RECT 1419.560 1700.000 1419.860 1700.340 ;
        RECT 1419.720 1684.350 1419.860 1700.000 ;
        RECT 1416.440 1684.030 1416.700 1684.350 ;
        RECT 1419.660 1684.030 1419.920 1684.350 ;
        RECT 1416.500 1677.290 1416.640 1684.030 ;
        RECT 1416.040 1677.150 1416.640 1677.290 ;
        RECT 1416.040 1349.110 1416.180 1677.150 ;
        RECT 1415.980 1348.790 1416.240 1349.110 ;
        RECT 2622.100 1348.790 2622.360 1349.110 ;
        RECT 2622.160 17.410 2622.300 1348.790 ;
        RECT 2622.160 17.270 2625.520 17.410 ;
        RECT 2625.380 2.400 2625.520 17.270 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1421.470 1683.920 1421.790 1683.980 ;
        RECT 1421.470 1683.780 1424.460 1683.920 ;
        RECT 1421.470 1683.720 1421.790 1683.780 ;
        RECT 1424.320 1683.580 1424.460 1683.780 ;
        RECT 1426.530 1683.580 1426.850 1683.640 ;
        RECT 1424.320 1683.440 1426.850 1683.580 ;
        RECT 1426.530 1683.380 1426.850 1683.440 ;
        RECT 1426.530 1341.880 1426.850 1341.940 ;
        RECT 2643.230 1341.880 2643.550 1341.940 ;
        RECT 1426.530 1341.740 2643.550 1341.880 ;
        RECT 1426.530 1341.680 1426.850 1341.740 ;
        RECT 2643.230 1341.680 2643.550 1341.740 ;
      LAYER via ;
        RECT 1421.500 1683.720 1421.760 1683.980 ;
        RECT 1426.560 1683.380 1426.820 1683.640 ;
        RECT 1426.560 1341.680 1426.820 1341.940 ;
        RECT 2643.260 1341.680 2643.520 1341.940 ;
      LAYER met2 ;
        RECT 1421.400 1700.340 1421.680 1704.000 ;
        RECT 1421.400 1700.000 1421.700 1700.340 ;
        RECT 1421.560 1684.010 1421.700 1700.000 ;
        RECT 1421.500 1683.690 1421.760 1684.010 ;
        RECT 1426.560 1683.350 1426.820 1683.670 ;
        RECT 1426.620 1341.970 1426.760 1683.350 ;
        RECT 1426.560 1341.650 1426.820 1341.970 ;
        RECT 2643.260 1341.650 2643.520 1341.970 ;
        RECT 2643.320 2.400 2643.460 1341.650 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1422.925 1442.025 1423.095 1490.475 ;
      LAYER mcon ;
        RECT 1422.925 1490.305 1423.095 1490.475 ;
      LAYER met1 ;
        RECT 1422.865 1490.460 1423.155 1490.505 ;
        RECT 1423.310 1490.460 1423.630 1490.520 ;
        RECT 1422.865 1490.320 1423.630 1490.460 ;
        RECT 1422.865 1490.275 1423.155 1490.320 ;
        RECT 1423.310 1490.260 1423.630 1490.320 ;
        RECT 1422.850 1442.180 1423.170 1442.240 ;
        RECT 1422.655 1442.040 1423.170 1442.180 ;
        RECT 1422.850 1441.980 1423.170 1442.040 ;
        RECT 1423.310 1335.080 1423.630 1335.140 ;
        RECT 2656.570 1335.080 2656.890 1335.140 ;
        RECT 1423.310 1334.940 2656.890 1335.080 ;
        RECT 1423.310 1334.880 1423.630 1334.940 ;
        RECT 2656.570 1334.880 2656.890 1334.940 ;
      LAYER via ;
        RECT 1423.340 1490.260 1423.600 1490.520 ;
        RECT 1422.880 1441.980 1423.140 1442.240 ;
        RECT 1423.340 1334.880 1423.600 1335.140 ;
        RECT 2656.600 1334.880 2656.860 1335.140 ;
      LAYER met2 ;
        RECT 1423.240 1700.410 1423.520 1704.000 ;
        RECT 1423.240 1700.270 1424.000 1700.410 ;
        RECT 1423.240 1700.000 1423.520 1700.270 ;
        RECT 1423.860 1632.410 1424.000 1700.270 ;
        RECT 1423.400 1632.270 1424.000 1632.410 ;
        RECT 1423.400 1490.550 1423.540 1632.270 ;
        RECT 1423.340 1490.230 1423.600 1490.550 ;
        RECT 1422.880 1441.950 1423.140 1442.270 ;
        RECT 1422.940 1414.810 1423.080 1441.950 ;
        RECT 1422.480 1414.670 1423.080 1414.810 ;
        RECT 1422.480 1414.130 1422.620 1414.670 ;
        RECT 1422.480 1413.990 1423.080 1414.130 ;
        RECT 1422.940 1366.530 1423.080 1413.990 ;
        RECT 1422.940 1366.390 1423.540 1366.530 ;
        RECT 1423.400 1335.170 1423.540 1366.390 ;
        RECT 1423.340 1334.850 1423.600 1335.170 ;
        RECT 2656.600 1334.850 2656.860 1335.170 ;
        RECT 2656.660 17.410 2656.800 1334.850 ;
        RECT 2656.660 17.270 2661.400 17.410 ;
        RECT 2661.260 2.400 2661.400 17.270 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1423.770 1631.900 1424.090 1631.960 ;
        RECT 1425.150 1631.900 1425.470 1631.960 ;
        RECT 1423.770 1631.760 1425.470 1631.900 ;
        RECT 1423.770 1631.700 1424.090 1631.760 ;
        RECT 1425.150 1631.700 1425.470 1631.760 ;
        RECT 1423.770 1328.280 1424.090 1328.340 ;
        RECT 2677.270 1328.280 2677.590 1328.340 ;
        RECT 1423.770 1328.140 2677.590 1328.280 ;
        RECT 1423.770 1328.080 1424.090 1328.140 ;
        RECT 2677.270 1328.080 2677.590 1328.140 ;
      LAYER via ;
        RECT 1423.800 1631.700 1424.060 1631.960 ;
        RECT 1425.180 1631.700 1425.440 1631.960 ;
        RECT 1423.800 1328.080 1424.060 1328.340 ;
        RECT 2677.300 1328.080 2677.560 1328.340 ;
      LAYER met2 ;
        RECT 1425.080 1700.340 1425.360 1704.000 ;
        RECT 1425.080 1700.000 1425.380 1700.340 ;
        RECT 1425.240 1631.990 1425.380 1700.000 ;
        RECT 1423.800 1631.670 1424.060 1631.990 ;
        RECT 1425.180 1631.670 1425.440 1631.990 ;
        RECT 1423.860 1328.370 1424.000 1631.670 ;
        RECT 1423.800 1328.050 1424.060 1328.370 ;
        RECT 2677.300 1328.050 2677.560 1328.370 ;
        RECT 2677.360 17.410 2677.500 1328.050 ;
        RECT 2677.360 17.270 2678.880 17.410 ;
        RECT 2678.740 2.400 2678.880 17.270 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1421.930 1685.960 1422.250 1686.020 ;
        RECT 1426.990 1685.960 1427.310 1686.020 ;
        RECT 1421.930 1685.820 1427.310 1685.960 ;
        RECT 1421.930 1685.760 1422.250 1685.820 ;
        RECT 1426.990 1685.760 1427.310 1685.820 ;
        RECT 1421.930 1631.560 1422.250 1631.620 ;
        RECT 1424.230 1631.560 1424.550 1631.620 ;
        RECT 1421.930 1631.420 1424.550 1631.560 ;
        RECT 1421.930 1631.360 1422.250 1631.420 ;
        RECT 1424.230 1631.360 1424.550 1631.420 ;
        RECT 1424.230 914.160 1424.550 914.220 ;
        RECT 2691.070 914.160 2691.390 914.220 ;
        RECT 1424.230 914.020 2691.390 914.160 ;
        RECT 1424.230 913.960 1424.550 914.020 ;
        RECT 2691.070 913.960 2691.390 914.020 ;
      LAYER via ;
        RECT 1421.960 1685.760 1422.220 1686.020 ;
        RECT 1427.020 1685.760 1427.280 1686.020 ;
        RECT 1421.960 1631.360 1422.220 1631.620 ;
        RECT 1424.260 1631.360 1424.520 1631.620 ;
        RECT 1424.260 913.960 1424.520 914.220 ;
        RECT 2691.100 913.960 2691.360 914.220 ;
      LAYER met2 ;
        RECT 1426.920 1700.340 1427.200 1704.000 ;
        RECT 1426.920 1700.000 1427.220 1700.340 ;
        RECT 1427.080 1686.050 1427.220 1700.000 ;
        RECT 1421.960 1685.730 1422.220 1686.050 ;
        RECT 1427.020 1685.730 1427.280 1686.050 ;
        RECT 1422.020 1631.650 1422.160 1685.730 ;
        RECT 1421.960 1631.330 1422.220 1631.650 ;
        RECT 1424.260 1631.330 1424.520 1631.650 ;
        RECT 1424.320 914.250 1424.460 1631.330 ;
        RECT 1424.260 913.930 1424.520 914.250 ;
        RECT 2691.100 913.930 2691.360 914.250 ;
        RECT 2691.160 17.410 2691.300 913.930 ;
        RECT 2691.160 17.270 2696.820 17.410 ;
        RECT 2696.680 2.400 2696.820 17.270 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1428.830 1452.380 1429.150 1452.440 ;
        RECT 2711.770 1452.380 2712.090 1452.440 ;
        RECT 1428.830 1452.240 2712.090 1452.380 ;
        RECT 1428.830 1452.180 1429.150 1452.240 ;
        RECT 2711.770 1452.180 2712.090 1452.240 ;
      LAYER via ;
        RECT 1428.860 1452.180 1429.120 1452.440 ;
        RECT 2711.800 1452.180 2712.060 1452.440 ;
      LAYER met2 ;
        RECT 1428.760 1700.340 1429.040 1704.000 ;
        RECT 1428.760 1700.000 1429.060 1700.340 ;
        RECT 1428.920 1452.470 1429.060 1700.000 ;
        RECT 1428.860 1452.150 1429.120 1452.470 ;
        RECT 2711.800 1452.150 2712.060 1452.470 ;
        RECT 2711.860 17.410 2712.000 1452.150 ;
        RECT 2711.860 17.270 2714.760 17.410 ;
        RECT 2714.620 2.400 2714.760 17.270 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1429.750 1314.340 1430.070 1314.400 ;
        RECT 2732.930 1314.340 2733.250 1314.400 ;
        RECT 1429.750 1314.200 2733.250 1314.340 ;
        RECT 1429.750 1314.140 1430.070 1314.200 ;
        RECT 2732.930 1314.140 2733.250 1314.200 ;
      LAYER via ;
        RECT 1429.780 1314.140 1430.040 1314.400 ;
        RECT 2732.960 1314.140 2733.220 1314.400 ;
      LAYER met2 ;
        RECT 1430.600 1700.340 1430.880 1704.000 ;
        RECT 1430.600 1700.000 1430.900 1700.340 ;
        RECT 1430.760 1677.970 1430.900 1700.000 ;
        RECT 1429.840 1677.830 1430.900 1677.970 ;
        RECT 1429.840 1314.430 1429.980 1677.830 ;
        RECT 1429.780 1314.110 1430.040 1314.430 ;
        RECT 2732.960 1314.110 2733.220 1314.430 ;
        RECT 2733.020 17.410 2733.160 1314.110 ;
        RECT 2732.560 17.270 2733.160 17.410 ;
        RECT 2732.560 2.400 2732.700 17.270 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1431.130 1684.260 1431.450 1684.320 ;
        RECT 1432.510 1684.260 1432.830 1684.320 ;
        RECT 1431.130 1684.120 1432.830 1684.260 ;
        RECT 1431.130 1684.060 1431.450 1684.120 ;
        RECT 1432.510 1684.060 1432.830 1684.120 ;
        RECT 1430.210 1307.540 1430.530 1307.600 ;
        RECT 2746.270 1307.540 2746.590 1307.600 ;
        RECT 1430.210 1307.400 2746.590 1307.540 ;
        RECT 1430.210 1307.340 1430.530 1307.400 ;
        RECT 2746.270 1307.340 2746.590 1307.400 ;
      LAYER via ;
        RECT 1431.160 1684.060 1431.420 1684.320 ;
        RECT 1432.540 1684.060 1432.800 1684.320 ;
        RECT 1430.240 1307.340 1430.500 1307.600 ;
        RECT 2746.300 1307.340 2746.560 1307.600 ;
      LAYER met2 ;
        RECT 1432.440 1700.340 1432.720 1704.000 ;
        RECT 1432.440 1700.000 1432.740 1700.340 ;
        RECT 1432.600 1684.350 1432.740 1700.000 ;
        RECT 1431.160 1684.030 1431.420 1684.350 ;
        RECT 1432.540 1684.030 1432.800 1684.350 ;
        RECT 1431.220 1677.290 1431.360 1684.030 ;
        RECT 1430.300 1677.150 1431.360 1677.290 ;
        RECT 1430.300 1307.630 1430.440 1677.150 ;
        RECT 1430.240 1307.310 1430.500 1307.630 ;
        RECT 2746.300 1307.310 2746.560 1307.630 ;
        RECT 2746.360 17.410 2746.500 1307.310 ;
        RECT 2746.360 17.270 2750.640 17.410 ;
        RECT 2750.500 2.400 2750.640 17.270 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1430.670 1676.780 1430.990 1676.840 ;
        RECT 1434.350 1676.780 1434.670 1676.840 ;
        RECT 1430.670 1676.640 1434.670 1676.780 ;
        RECT 1430.670 1676.580 1430.990 1676.640 ;
        RECT 1434.350 1676.580 1434.670 1676.640 ;
        RECT 1430.670 1300.740 1430.990 1300.800 ;
        RECT 2766.970 1300.740 2767.290 1300.800 ;
        RECT 1430.670 1300.600 2767.290 1300.740 ;
        RECT 1430.670 1300.540 1430.990 1300.600 ;
        RECT 2766.970 1300.540 2767.290 1300.600 ;
      LAYER via ;
        RECT 1430.700 1676.580 1430.960 1676.840 ;
        RECT 1434.380 1676.580 1434.640 1676.840 ;
        RECT 1430.700 1300.540 1430.960 1300.800 ;
        RECT 2767.000 1300.540 2767.260 1300.800 ;
      LAYER met2 ;
        RECT 1434.280 1700.340 1434.560 1704.000 ;
        RECT 1434.280 1700.000 1434.580 1700.340 ;
        RECT 1434.440 1676.870 1434.580 1700.000 ;
        RECT 1430.700 1676.550 1430.960 1676.870 ;
        RECT 1434.380 1676.550 1434.640 1676.870 ;
        RECT 1430.760 1300.830 1430.900 1676.550 ;
        RECT 1430.700 1300.510 1430.960 1300.830 ;
        RECT 2767.000 1300.510 2767.260 1300.830 ;
        RECT 2767.060 17.410 2767.200 1300.510 ;
        RECT 2767.060 17.270 2768.120 17.410 ;
        RECT 2767.980 2.400 2768.120 17.270 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 840.950 38.320 841.270 38.380 ;
        RECT 1237.470 38.320 1237.790 38.380 ;
        RECT 840.950 38.180 1237.790 38.320 ;
        RECT 840.950 38.120 841.270 38.180 ;
        RECT 1237.470 38.120 1237.790 38.180 ;
      LAYER via ;
        RECT 840.980 38.120 841.240 38.380 ;
        RECT 1237.500 38.120 1237.760 38.380 ;
      LAYER met2 ;
        RECT 1236.020 1700.340 1236.300 1704.000 ;
        RECT 1236.020 1700.000 1236.320 1700.340 ;
        RECT 1236.180 1667.770 1236.320 1700.000 ;
        RECT 1236.180 1667.630 1237.700 1667.770 ;
        RECT 1237.560 38.410 1237.700 1667.630 ;
        RECT 840.980 38.090 841.240 38.410 ;
        RECT 1237.500 38.090 1237.760 38.410 ;
        RECT 841.040 2.400 841.180 38.090 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1441.785 1445.425 1441.955 1490.475 ;
      LAYER mcon ;
        RECT 1441.785 1490.305 1441.955 1490.475 ;
      LAYER met1 ;
        RECT 1437.110 1656.380 1437.430 1656.440 ;
        RECT 1437.110 1656.240 1440.100 1656.380 ;
        RECT 1437.110 1656.180 1437.430 1656.240 ;
        RECT 1439.960 1656.100 1440.100 1656.240 ;
        RECT 1439.870 1655.840 1440.190 1656.100 ;
        RECT 1441.710 1490.460 1442.030 1490.520 ;
        RECT 1441.515 1490.320 1442.030 1490.460 ;
        RECT 1441.710 1490.260 1442.030 1490.320 ;
        RECT 1441.725 1445.580 1442.015 1445.625 ;
        RECT 2780.770 1445.580 2781.090 1445.640 ;
        RECT 1441.725 1445.440 2781.090 1445.580 ;
        RECT 1441.725 1445.395 1442.015 1445.440 ;
        RECT 2780.770 1445.380 2781.090 1445.440 ;
      LAYER via ;
        RECT 1437.140 1656.180 1437.400 1656.440 ;
        RECT 1439.900 1655.840 1440.160 1656.100 ;
        RECT 1441.740 1490.260 1442.000 1490.520 ;
        RECT 2780.800 1445.380 2781.060 1445.640 ;
      LAYER met2 ;
        RECT 1436.120 1700.340 1436.400 1704.000 ;
        RECT 1436.120 1700.000 1436.420 1700.340 ;
        RECT 1436.280 1684.770 1436.420 1700.000 ;
        RECT 1436.280 1684.630 1437.340 1684.770 ;
        RECT 1437.200 1656.470 1437.340 1684.630 ;
        RECT 1437.140 1656.150 1437.400 1656.470 ;
        RECT 1439.900 1655.810 1440.160 1656.130 ;
        RECT 1439.960 1624.250 1440.100 1655.810 ;
        RECT 1439.960 1624.110 1441.020 1624.250 ;
        RECT 1440.880 1569.850 1441.020 1624.110 ;
        RECT 1440.880 1569.710 1441.940 1569.850 ;
        RECT 1441.800 1490.550 1441.940 1569.710 ;
        RECT 1441.740 1490.230 1442.000 1490.550 ;
        RECT 2780.800 1445.350 2781.060 1445.670 ;
        RECT 2780.860 18.090 2781.000 1445.350 ;
        RECT 2780.860 17.950 2786.060 18.090 ;
        RECT 2785.920 2.400 2786.060 17.950 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1436.190 1683.920 1436.510 1683.980 ;
        RECT 1438.030 1683.920 1438.350 1683.980 ;
        RECT 1436.190 1683.780 1438.350 1683.920 ;
        RECT 1436.190 1683.720 1436.510 1683.780 ;
        RECT 1438.030 1683.720 1438.350 1683.780 ;
        RECT 1436.190 1293.600 1436.510 1293.660 ;
        RECT 2801.470 1293.600 2801.790 1293.660 ;
        RECT 1436.190 1293.460 2801.790 1293.600 ;
        RECT 1436.190 1293.400 1436.510 1293.460 ;
        RECT 2801.470 1293.400 2801.790 1293.460 ;
      LAYER via ;
        RECT 1436.220 1683.720 1436.480 1683.980 ;
        RECT 1438.060 1683.720 1438.320 1683.980 ;
        RECT 1436.220 1293.400 1436.480 1293.660 ;
        RECT 2801.500 1293.400 2801.760 1293.660 ;
      LAYER met2 ;
        RECT 1437.960 1700.340 1438.240 1704.000 ;
        RECT 1437.960 1700.000 1438.260 1700.340 ;
        RECT 1438.120 1684.010 1438.260 1700.000 ;
        RECT 1436.220 1683.690 1436.480 1684.010 ;
        RECT 1438.060 1683.690 1438.320 1684.010 ;
        RECT 1436.280 1293.690 1436.420 1683.690 ;
        RECT 1436.220 1293.370 1436.480 1293.690 ;
        RECT 2801.500 1293.370 2801.760 1293.690 ;
        RECT 2801.560 17.410 2801.700 1293.370 ;
        RECT 2801.560 17.270 2804.000 17.410 ;
        RECT 2803.860 2.400 2804.000 17.270 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1436.650 1684.260 1436.970 1684.320 ;
        RECT 1439.870 1684.260 1440.190 1684.320 ;
        RECT 1436.650 1684.120 1440.190 1684.260 ;
        RECT 1436.650 1684.060 1436.970 1684.120 ;
        RECT 1439.870 1684.060 1440.190 1684.120 ;
        RECT 1436.650 1286.800 1436.970 1286.860 ;
        RECT 2815.730 1286.800 2816.050 1286.860 ;
        RECT 1436.650 1286.660 2816.050 1286.800 ;
        RECT 1436.650 1286.600 1436.970 1286.660 ;
        RECT 2815.730 1286.600 2816.050 1286.660 ;
        RECT 2815.730 18.260 2816.050 18.320 ;
        RECT 2821.710 18.260 2822.030 18.320 ;
        RECT 2815.730 18.120 2822.030 18.260 ;
        RECT 2815.730 18.060 2816.050 18.120 ;
        RECT 2821.710 18.060 2822.030 18.120 ;
      LAYER via ;
        RECT 1436.680 1684.060 1436.940 1684.320 ;
        RECT 1439.900 1684.060 1440.160 1684.320 ;
        RECT 1436.680 1286.600 1436.940 1286.860 ;
        RECT 2815.760 1286.600 2816.020 1286.860 ;
        RECT 2815.760 18.060 2816.020 18.320 ;
        RECT 2821.740 18.060 2822.000 18.320 ;
      LAYER met2 ;
        RECT 1439.800 1700.340 1440.080 1704.000 ;
        RECT 1439.800 1700.000 1440.100 1700.340 ;
        RECT 1439.960 1684.350 1440.100 1700.000 ;
        RECT 1436.680 1684.030 1436.940 1684.350 ;
        RECT 1439.900 1684.030 1440.160 1684.350 ;
        RECT 1436.740 1286.890 1436.880 1684.030 ;
        RECT 1436.680 1286.570 1436.940 1286.890 ;
        RECT 2815.760 1286.570 2816.020 1286.890 ;
        RECT 2815.820 18.350 2815.960 1286.570 ;
        RECT 2815.760 18.030 2816.020 18.350 ;
        RECT 2821.740 18.030 2822.000 18.350 ;
        RECT 2821.800 2.400 2821.940 18.030 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1438.030 1631.560 1438.350 1631.620 ;
        RECT 1441.710 1631.560 1442.030 1631.620 ;
        RECT 1438.030 1631.420 1442.030 1631.560 ;
        RECT 1438.030 1631.360 1438.350 1631.420 ;
        RECT 1441.710 1631.360 1442.030 1631.420 ;
        RECT 1438.030 141.340 1438.350 141.400 ;
        RECT 2835.970 141.340 2836.290 141.400 ;
        RECT 1438.030 141.200 2836.290 141.340 ;
        RECT 1438.030 141.140 1438.350 141.200 ;
        RECT 2835.970 141.140 2836.290 141.200 ;
      LAYER via ;
        RECT 1438.060 1631.360 1438.320 1631.620 ;
        RECT 1441.740 1631.360 1442.000 1631.620 ;
        RECT 1438.060 141.140 1438.320 141.400 ;
        RECT 2836.000 141.140 2836.260 141.400 ;
      LAYER met2 ;
        RECT 1441.640 1700.340 1441.920 1704.000 ;
        RECT 1441.640 1700.000 1441.940 1700.340 ;
        RECT 1441.800 1631.650 1441.940 1700.000 ;
        RECT 1438.060 1631.330 1438.320 1631.650 ;
        RECT 1441.740 1631.330 1442.000 1631.650 ;
        RECT 1438.120 141.430 1438.260 1631.330 ;
        RECT 1438.060 141.110 1438.320 141.430 ;
        RECT 2836.000 141.110 2836.260 141.430 ;
        RECT 2836.060 16.730 2836.200 141.110 ;
        RECT 2836.060 16.590 2839.420 16.730 ;
        RECT 2839.280 2.400 2839.420 16.590 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1443.550 1487.060 1443.870 1487.120 ;
        RECT 2852.990 1487.060 2853.310 1487.120 ;
        RECT 1443.550 1486.920 2853.310 1487.060 ;
        RECT 1443.550 1486.860 1443.870 1486.920 ;
        RECT 2852.990 1486.860 2853.310 1486.920 ;
        RECT 2852.990 17.920 2853.310 17.980 ;
        RECT 2857.130 17.920 2857.450 17.980 ;
        RECT 2852.990 17.780 2857.450 17.920 ;
        RECT 2852.990 17.720 2853.310 17.780 ;
        RECT 2857.130 17.720 2857.450 17.780 ;
      LAYER via ;
        RECT 1443.580 1486.860 1443.840 1487.120 ;
        RECT 2853.020 1486.860 2853.280 1487.120 ;
        RECT 2853.020 17.720 2853.280 17.980 ;
        RECT 2857.160 17.720 2857.420 17.980 ;
      LAYER met2 ;
        RECT 1443.480 1700.340 1443.760 1704.000 ;
        RECT 1443.480 1700.000 1443.780 1700.340 ;
        RECT 1443.640 1487.150 1443.780 1700.000 ;
        RECT 1443.580 1486.830 1443.840 1487.150 ;
        RECT 2853.020 1486.830 2853.280 1487.150 ;
        RECT 2853.080 18.010 2853.220 1486.830 ;
        RECT 2853.020 17.690 2853.280 18.010 ;
        RECT 2857.160 17.690 2857.420 18.010 ;
        RECT 2857.220 2.400 2857.360 17.690 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2838.805 16.745 2838.975 17.935 ;
      LAYER mcon ;
        RECT 2838.805 17.765 2838.975 17.935 ;
      LAYER met1 ;
        RECT 1445.390 1608.440 1445.710 1608.500 ;
        RECT 1445.020 1608.300 1445.710 1608.440 ;
        RECT 1445.020 1607.820 1445.160 1608.300 ;
        RECT 1445.390 1608.240 1445.710 1608.300 ;
        RECT 1444.930 1607.560 1445.250 1607.820 ;
        RECT 1444.930 1480.260 1445.250 1480.320 ;
        RECT 2411.390 1480.260 2411.710 1480.320 ;
        RECT 1444.930 1480.120 2411.710 1480.260 ;
        RECT 1444.930 1480.060 1445.250 1480.120 ;
        RECT 2411.390 1480.060 2411.710 1480.120 ;
        RECT 2411.390 17.920 2411.710 17.980 ;
        RECT 2838.745 17.920 2839.035 17.965 ;
        RECT 2411.390 17.780 2839.035 17.920 ;
        RECT 2411.390 17.720 2411.710 17.780 ;
        RECT 2838.745 17.735 2839.035 17.780 ;
        RECT 2838.745 16.900 2839.035 16.945 ;
        RECT 2875.070 16.900 2875.390 16.960 ;
        RECT 2838.745 16.760 2875.390 16.900 ;
        RECT 2838.745 16.715 2839.035 16.760 ;
        RECT 2875.070 16.700 2875.390 16.760 ;
      LAYER via ;
        RECT 1445.420 1608.240 1445.680 1608.500 ;
        RECT 1444.960 1607.560 1445.220 1607.820 ;
        RECT 1444.960 1480.060 1445.220 1480.320 ;
        RECT 2411.420 1480.060 2411.680 1480.320 ;
        RECT 2411.420 17.720 2411.680 17.980 ;
        RECT 2875.100 16.700 2875.360 16.960 ;
      LAYER met2 ;
        RECT 1445.320 1700.340 1445.600 1704.000 ;
        RECT 1445.320 1700.000 1445.620 1700.340 ;
        RECT 1445.480 1608.530 1445.620 1700.000 ;
        RECT 1445.420 1608.210 1445.680 1608.530 ;
        RECT 1444.960 1607.530 1445.220 1607.850 ;
        RECT 1445.020 1480.350 1445.160 1607.530 ;
        RECT 1444.960 1480.030 1445.220 1480.350 ;
        RECT 2411.420 1480.030 2411.680 1480.350 ;
        RECT 2411.480 18.010 2411.620 1480.030 ;
        RECT 2411.420 17.690 2411.680 18.010 ;
        RECT 2875.100 16.670 2875.360 16.990 ;
        RECT 2875.160 2.400 2875.300 16.670 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1445.925 1594.005 1446.095 1617.975 ;
        RECT 1445.465 1442.025 1445.635 1490.475 ;
      LAYER mcon ;
        RECT 1445.925 1617.805 1446.095 1617.975 ;
        RECT 1445.465 1490.305 1445.635 1490.475 ;
      LAYER met1 ;
        RECT 1445.850 1617.960 1446.170 1618.020 ;
        RECT 1445.655 1617.820 1446.170 1617.960 ;
        RECT 1445.850 1617.760 1446.170 1617.820 ;
        RECT 1445.865 1594.160 1446.155 1594.205 ;
        RECT 1446.310 1594.160 1446.630 1594.220 ;
        RECT 1445.865 1594.020 1446.630 1594.160 ;
        RECT 1445.865 1593.975 1446.155 1594.020 ;
        RECT 1446.310 1593.960 1446.630 1594.020 ;
        RECT 1445.405 1490.460 1445.695 1490.505 ;
        RECT 1446.310 1490.460 1446.630 1490.520 ;
        RECT 1445.405 1490.320 1446.630 1490.460 ;
        RECT 1445.405 1490.275 1445.695 1490.320 ;
        RECT 1446.310 1490.260 1446.630 1490.320 ;
        RECT 1445.390 1442.180 1445.710 1442.240 ;
        RECT 1445.195 1442.040 1445.710 1442.180 ;
        RECT 1445.390 1441.980 1445.710 1442.040 ;
        RECT 1444.470 1321.140 1444.790 1321.200 ;
        RECT 2376.890 1321.140 2377.210 1321.200 ;
        RECT 1444.470 1321.000 2377.210 1321.140 ;
        RECT 1444.470 1320.940 1444.790 1321.000 ;
        RECT 2376.890 1320.940 2377.210 1321.000 ;
        RECT 2376.890 17.580 2377.210 17.640 ;
        RECT 2893.010 17.580 2893.330 17.640 ;
        RECT 2376.890 17.440 2893.330 17.580 ;
        RECT 2376.890 17.380 2377.210 17.440 ;
        RECT 2893.010 17.380 2893.330 17.440 ;
      LAYER via ;
        RECT 1445.880 1617.760 1446.140 1618.020 ;
        RECT 1446.340 1593.960 1446.600 1594.220 ;
        RECT 1446.340 1490.260 1446.600 1490.520 ;
        RECT 1445.420 1441.980 1445.680 1442.240 ;
        RECT 1444.500 1320.940 1444.760 1321.200 ;
        RECT 2376.920 1320.940 2377.180 1321.200 ;
        RECT 2376.920 17.380 2377.180 17.640 ;
        RECT 2893.040 17.380 2893.300 17.640 ;
      LAYER met2 ;
        RECT 1447.160 1700.340 1447.440 1704.000 ;
        RECT 1447.160 1700.000 1447.460 1700.340 ;
        RECT 1447.320 1677.970 1447.460 1700.000 ;
        RECT 1445.940 1677.830 1447.460 1677.970 ;
        RECT 1445.940 1618.050 1446.080 1677.830 ;
        RECT 1445.880 1617.730 1446.140 1618.050 ;
        RECT 1446.340 1593.930 1446.600 1594.250 ;
        RECT 1446.400 1490.550 1446.540 1593.930 ;
        RECT 1446.340 1490.230 1446.600 1490.550 ;
        RECT 1445.420 1441.950 1445.680 1442.270 ;
        RECT 1445.480 1414.810 1445.620 1441.950 ;
        RECT 1444.560 1414.670 1445.620 1414.810 ;
        RECT 1444.560 1321.230 1444.700 1414.670 ;
        RECT 1444.500 1320.910 1444.760 1321.230 ;
        RECT 2376.920 1320.910 2377.180 1321.230 ;
        RECT 2376.980 17.670 2377.120 1320.910 ;
        RECT 2376.920 17.350 2377.180 17.670 ;
        RECT 2893.040 17.350 2893.300 17.670 ;
        RECT 2893.100 2.400 2893.240 17.350 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1455.510 1280.000 1455.830 1280.060 ;
        RECT 2356.190 1280.000 2356.510 1280.060 ;
        RECT 1455.510 1279.860 2356.510 1280.000 ;
        RECT 1455.510 1279.800 1455.830 1279.860 ;
        RECT 2356.190 1279.800 2356.510 1279.860 ;
        RECT 2356.190 17.240 2356.510 17.300 ;
        RECT 2910.950 17.240 2911.270 17.300 ;
        RECT 2356.190 17.100 2911.270 17.240 ;
        RECT 2356.190 17.040 2356.510 17.100 ;
        RECT 2910.950 17.040 2911.270 17.100 ;
      LAYER via ;
        RECT 1455.540 1279.800 1455.800 1280.060 ;
        RECT 2356.220 1279.800 2356.480 1280.060 ;
        RECT 2356.220 17.040 2356.480 17.300 ;
        RECT 2910.980 17.040 2911.240 17.300 ;
      LAYER met2 ;
        RECT 1449.000 1700.340 1449.280 1704.000 ;
        RECT 1449.000 1700.000 1449.300 1700.340 ;
        RECT 1449.160 1689.645 1449.300 1700.000 ;
        RECT 1449.090 1689.275 1449.370 1689.645 ;
        RECT 1455.530 1689.275 1455.810 1689.645 ;
        RECT 1455.600 1280.090 1455.740 1689.275 ;
        RECT 1455.540 1279.770 1455.800 1280.090 ;
        RECT 2356.220 1279.770 2356.480 1280.090 ;
        RECT 2356.280 17.330 2356.420 1279.770 ;
        RECT 2356.220 17.010 2356.480 17.330 ;
        RECT 2910.980 17.010 2911.240 17.330 ;
        RECT 2911.040 2.400 2911.180 17.010 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
      LAYER via2 ;
        RECT 1449.090 1689.320 1449.370 1689.600 ;
        RECT 1455.530 1689.320 1455.810 1689.600 ;
      LAYER met3 ;
        RECT 1449.065 1689.610 1449.395 1689.625 ;
        RECT 1455.505 1689.610 1455.835 1689.625 ;
        RECT 1449.065 1689.310 1455.835 1689.610 ;
        RECT 1449.065 1689.295 1449.395 1689.310 ;
        RECT 1455.505 1689.295 1455.835 1689.310 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1237.930 1678.140 1238.250 1678.200 ;
        RECT 1239.310 1678.140 1239.630 1678.200 ;
        RECT 1237.930 1678.000 1239.630 1678.140 ;
        RECT 1237.930 1677.940 1238.250 1678.000 ;
        RECT 1239.310 1677.940 1239.630 1678.000 ;
        RECT 858.890 38.660 859.210 38.720 ;
        RECT 1239.310 38.660 1239.630 38.720 ;
        RECT 858.890 38.520 1239.630 38.660 ;
        RECT 858.890 38.460 859.210 38.520 ;
        RECT 1239.310 38.460 1239.630 38.520 ;
      LAYER via ;
        RECT 1237.960 1677.940 1238.220 1678.200 ;
        RECT 1239.340 1677.940 1239.600 1678.200 ;
        RECT 858.920 38.460 859.180 38.720 ;
        RECT 1239.340 38.460 1239.600 38.720 ;
      LAYER met2 ;
        RECT 1237.860 1700.340 1238.140 1704.000 ;
        RECT 1237.860 1700.000 1238.160 1700.340 ;
        RECT 1238.020 1678.230 1238.160 1700.000 ;
        RECT 1237.960 1677.910 1238.220 1678.230 ;
        RECT 1239.340 1677.910 1239.600 1678.230 ;
        RECT 1239.400 38.750 1239.540 1677.910 ;
        RECT 858.920 38.430 859.180 38.750 ;
        RECT 1239.340 38.430 1239.600 38.750 ;
        RECT 858.980 2.400 859.120 38.430 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1236.550 1667.260 1236.870 1667.320 ;
        RECT 1239.770 1667.260 1240.090 1667.320 ;
        RECT 1236.550 1667.120 1240.090 1667.260 ;
        RECT 1236.550 1667.060 1236.870 1667.120 ;
        RECT 1239.770 1667.060 1240.090 1667.120 ;
        RECT 876.830 39.000 877.150 39.060 ;
        RECT 1236.550 39.000 1236.870 39.060 ;
        RECT 876.830 38.860 1236.870 39.000 ;
        RECT 876.830 38.800 877.150 38.860 ;
        RECT 1236.550 38.800 1236.870 38.860 ;
      LAYER via ;
        RECT 1236.580 1667.060 1236.840 1667.320 ;
        RECT 1239.800 1667.060 1240.060 1667.320 ;
        RECT 876.860 38.800 877.120 39.060 ;
        RECT 1236.580 38.800 1236.840 39.060 ;
      LAYER met2 ;
        RECT 1239.700 1700.340 1239.980 1704.000 ;
        RECT 1239.700 1700.000 1240.000 1700.340 ;
        RECT 1239.860 1667.350 1240.000 1700.000 ;
        RECT 1236.580 1667.030 1236.840 1667.350 ;
        RECT 1239.800 1667.030 1240.060 1667.350 ;
        RECT 1236.640 39.090 1236.780 1667.030 ;
        RECT 876.860 38.770 877.120 39.090 ;
        RECT 1236.580 38.770 1236.840 39.090 ;
        RECT 876.920 2.400 877.060 38.770 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1237.010 1666.920 1237.330 1666.980 ;
        RECT 1241.610 1666.920 1241.930 1666.980 ;
        RECT 1237.010 1666.780 1241.930 1666.920 ;
        RECT 1237.010 1666.720 1237.330 1666.780 ;
        RECT 1241.610 1666.720 1241.930 1666.780 ;
        RECT 894.770 39.340 895.090 39.400 ;
        RECT 1237.010 39.340 1237.330 39.400 ;
        RECT 894.770 39.200 1237.330 39.340 ;
        RECT 894.770 39.140 895.090 39.200 ;
        RECT 1237.010 39.140 1237.330 39.200 ;
      LAYER via ;
        RECT 1237.040 1666.720 1237.300 1666.980 ;
        RECT 1241.640 1666.720 1241.900 1666.980 ;
        RECT 894.800 39.140 895.060 39.400 ;
        RECT 1237.040 39.140 1237.300 39.400 ;
      LAYER met2 ;
        RECT 1241.540 1700.340 1241.820 1704.000 ;
        RECT 1241.540 1700.000 1241.840 1700.340 ;
        RECT 1241.700 1667.010 1241.840 1700.000 ;
        RECT 1237.040 1666.690 1237.300 1667.010 ;
        RECT 1241.640 1666.690 1241.900 1667.010 ;
        RECT 1237.100 39.430 1237.240 1666.690 ;
        RECT 894.800 39.110 895.060 39.430 ;
        RECT 1237.040 39.110 1237.300 39.430 ;
        RECT 894.860 2.400 895.000 39.110 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 912.710 39.680 913.030 39.740 ;
        RECT 1243.910 39.680 1244.230 39.740 ;
        RECT 912.710 39.540 1244.230 39.680 ;
        RECT 912.710 39.480 913.030 39.540 ;
        RECT 1243.910 39.480 1244.230 39.540 ;
      LAYER via ;
        RECT 912.740 39.480 913.000 39.740 ;
        RECT 1243.940 39.480 1244.200 39.740 ;
      LAYER met2 ;
        RECT 1243.380 1700.340 1243.660 1704.000 ;
        RECT 1243.380 1700.000 1243.680 1700.340 ;
        RECT 1243.540 1677.970 1243.680 1700.000 ;
        RECT 1243.540 1677.830 1244.140 1677.970 ;
        RECT 1244.000 39.770 1244.140 1677.830 ;
        RECT 912.740 39.450 913.000 39.770 ;
        RECT 1243.940 39.450 1244.200 39.770 ;
        RECT 912.800 2.400 912.940 39.450 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1243.450 1677.460 1243.770 1677.520 ;
        RECT 1245.290 1677.460 1245.610 1677.520 ;
        RECT 1243.450 1677.320 1245.610 1677.460 ;
        RECT 1243.450 1677.260 1243.770 1677.320 ;
        RECT 1245.290 1677.260 1245.610 1677.320 ;
        RECT 930.190 40.020 930.510 40.080 ;
        RECT 1243.450 40.020 1243.770 40.080 ;
        RECT 930.190 39.880 1243.770 40.020 ;
        RECT 930.190 39.820 930.510 39.880 ;
        RECT 1243.450 39.820 1243.770 39.880 ;
      LAYER via ;
        RECT 1243.480 1677.260 1243.740 1677.520 ;
        RECT 1245.320 1677.260 1245.580 1677.520 ;
        RECT 930.220 39.820 930.480 40.080 ;
        RECT 1243.480 39.820 1243.740 40.080 ;
      LAYER met2 ;
        RECT 1245.220 1700.340 1245.500 1704.000 ;
        RECT 1245.220 1700.000 1245.520 1700.340 ;
        RECT 1245.380 1677.550 1245.520 1700.000 ;
        RECT 1243.480 1677.230 1243.740 1677.550 ;
        RECT 1245.320 1677.230 1245.580 1677.550 ;
        RECT 1243.540 40.110 1243.680 1677.230 ;
        RECT 930.220 39.790 930.480 40.110 ;
        RECT 1243.480 39.790 1243.740 40.110 ;
        RECT 930.280 2.400 930.420 39.790 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 948.130 40.360 948.450 40.420 ;
        RECT 1247.130 40.360 1247.450 40.420 ;
        RECT 948.130 40.220 1247.450 40.360 ;
        RECT 948.130 40.160 948.450 40.220 ;
        RECT 1247.130 40.160 1247.450 40.220 ;
      LAYER via ;
        RECT 948.160 40.160 948.420 40.420 ;
        RECT 1247.160 40.160 1247.420 40.420 ;
      LAYER met2 ;
        RECT 1247.060 1700.340 1247.340 1704.000 ;
        RECT 1247.060 1700.000 1247.360 1700.340 ;
        RECT 1247.220 40.450 1247.360 1700.000 ;
        RECT 948.160 40.130 948.420 40.450 ;
        RECT 1247.160 40.130 1247.420 40.450 ;
        RECT 948.220 2.400 948.360 40.130 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 966.070 40.700 966.390 40.760 ;
        RECT 1249.430 40.700 1249.750 40.760 ;
        RECT 966.070 40.560 1249.750 40.700 ;
        RECT 966.070 40.500 966.390 40.560 ;
        RECT 1249.430 40.500 1249.750 40.560 ;
      LAYER via ;
        RECT 966.100 40.500 966.360 40.760 ;
        RECT 1249.460 40.500 1249.720 40.760 ;
      LAYER met2 ;
        RECT 1248.900 1700.340 1249.180 1704.000 ;
        RECT 1248.900 1700.000 1249.200 1700.340 ;
        RECT 1249.060 1677.970 1249.200 1700.000 ;
        RECT 1249.060 1677.830 1249.660 1677.970 ;
        RECT 1249.520 40.790 1249.660 1677.830 ;
        RECT 966.100 40.470 966.360 40.790 ;
        RECT 1249.460 40.470 1249.720 40.790 ;
        RECT 966.160 2.400 966.300 40.470 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 984.010 41.040 984.330 41.100 ;
        RECT 1250.810 41.040 1251.130 41.100 ;
        RECT 984.010 40.900 1251.130 41.040 ;
        RECT 984.010 40.840 984.330 40.900 ;
        RECT 1250.810 40.840 1251.130 40.900 ;
      LAYER via ;
        RECT 984.040 40.840 984.300 41.100 ;
        RECT 1250.840 40.840 1251.100 41.100 ;
      LAYER met2 ;
        RECT 1250.740 1700.340 1251.020 1704.000 ;
        RECT 1250.740 1700.000 1251.040 1700.340 ;
        RECT 1250.900 41.130 1251.040 1700.000 ;
        RECT 984.040 40.810 984.300 41.130 ;
        RECT 1250.840 40.810 1251.100 41.130 ;
        RECT 984.100 2.400 984.240 40.810 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1217.690 1463.260 1218.010 1463.320 ;
        RECT 1216.860 1463.120 1218.010 1463.260 ;
        RECT 1216.860 1462.980 1217.000 1463.120 ;
        RECT 1217.690 1463.060 1218.010 1463.120 ;
        RECT 1216.770 1462.720 1217.090 1462.980 ;
        RECT 1216.770 1172.900 1217.090 1172.960 ;
        RECT 1217.690 1172.900 1218.010 1172.960 ;
        RECT 1216.770 1172.760 1218.010 1172.900 ;
        RECT 1216.770 1172.700 1217.090 1172.760 ;
        RECT 1217.690 1172.700 1218.010 1172.760 ;
        RECT 1217.690 1077.020 1218.010 1077.080 ;
        RECT 1216.860 1076.880 1218.010 1077.020 ;
        RECT 1216.860 1076.740 1217.000 1076.880 ;
        RECT 1217.690 1076.820 1218.010 1076.880 ;
        RECT 1216.770 1076.480 1217.090 1076.740 ;
        RECT 1216.770 496.640 1217.090 496.700 ;
        RECT 1217.690 496.640 1218.010 496.700 ;
        RECT 1216.770 496.500 1218.010 496.640 ;
        RECT 1216.770 496.440 1217.090 496.500 ;
        RECT 1217.690 496.440 1218.010 496.500 ;
        RECT 1216.770 352.140 1217.090 352.200 ;
        RECT 1217.690 352.140 1218.010 352.200 ;
        RECT 1216.770 352.000 1218.010 352.140 ;
        RECT 1216.770 351.940 1217.090 352.000 ;
        RECT 1217.690 351.940 1218.010 352.000 ;
        RECT 662.930 37.980 663.250 38.040 ;
        RECT 1216.770 37.980 1217.090 38.040 ;
        RECT 662.930 37.840 1217.090 37.980 ;
        RECT 662.930 37.780 663.250 37.840 ;
        RECT 1216.770 37.780 1217.090 37.840 ;
      LAYER via ;
        RECT 1217.720 1463.060 1217.980 1463.320 ;
        RECT 1216.800 1462.720 1217.060 1462.980 ;
        RECT 1216.800 1172.700 1217.060 1172.960 ;
        RECT 1217.720 1172.700 1217.980 1172.960 ;
        RECT 1217.720 1076.820 1217.980 1077.080 ;
        RECT 1216.800 1076.480 1217.060 1076.740 ;
        RECT 1216.800 496.440 1217.060 496.700 ;
        RECT 1217.720 496.440 1217.980 496.700 ;
        RECT 1216.800 351.940 1217.060 352.200 ;
        RECT 1217.720 351.940 1217.980 352.200 ;
        RECT 662.960 37.780 663.220 38.040 ;
        RECT 1216.800 37.780 1217.060 38.040 ;
      LAYER met2 ;
        RECT 1217.620 1700.340 1217.900 1704.000 ;
        RECT 1217.620 1700.000 1217.920 1700.340 ;
        RECT 1217.780 1463.350 1217.920 1700.000 ;
        RECT 1217.720 1463.030 1217.980 1463.350 ;
        RECT 1216.800 1462.690 1217.060 1463.010 ;
        RECT 1216.860 1172.990 1217.000 1462.690 ;
        RECT 1216.800 1172.670 1217.060 1172.990 ;
        RECT 1217.720 1172.670 1217.980 1172.990 ;
        RECT 1217.780 1077.110 1217.920 1172.670 ;
        RECT 1217.720 1076.790 1217.980 1077.110 ;
        RECT 1216.800 1076.450 1217.060 1076.770 ;
        RECT 1216.860 496.730 1217.000 1076.450 ;
        RECT 1216.800 496.410 1217.060 496.730 ;
        RECT 1217.720 496.410 1217.980 496.730 ;
        RECT 1217.780 352.230 1217.920 496.410 ;
        RECT 1216.800 351.910 1217.060 352.230 ;
        RECT 1217.720 351.910 1217.980 352.230 ;
        RECT 1216.860 38.070 1217.000 351.910 ;
        RECT 662.960 37.750 663.220 38.070 ;
        RECT 1216.800 37.750 1217.060 38.070 ;
        RECT 663.020 2.400 663.160 37.750 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1252.725 1642.285 1252.895 1666.595 ;
        RECT 1253.645 1268.965 1253.815 1304.155 ;
        RECT 1252.725 641.325 1252.895 703.715 ;
        RECT 1253.185 510.765 1253.355 558.875 ;
        RECT 1253.645 341.445 1253.815 414.035 ;
        RECT 1252.265 48.365 1252.435 96.475 ;
      LAYER mcon ;
        RECT 1252.725 1666.425 1252.895 1666.595 ;
        RECT 1253.645 1303.985 1253.815 1304.155 ;
        RECT 1252.725 703.545 1252.895 703.715 ;
        RECT 1253.185 558.705 1253.355 558.875 ;
        RECT 1253.645 413.865 1253.815 414.035 ;
        RECT 1252.265 96.305 1252.435 96.475 ;
      LAYER met1 ;
        RECT 1252.650 1666.580 1252.970 1666.640 ;
        RECT 1252.455 1666.440 1252.970 1666.580 ;
        RECT 1252.650 1666.380 1252.970 1666.440 ;
        RECT 1252.665 1642.440 1252.955 1642.485 ;
        RECT 1253.110 1642.440 1253.430 1642.500 ;
        RECT 1252.665 1642.300 1253.430 1642.440 ;
        RECT 1252.665 1642.255 1252.955 1642.300 ;
        RECT 1253.110 1642.240 1253.430 1642.300 ;
        RECT 1252.650 1401.040 1252.970 1401.100 ;
        RECT 1253.570 1401.040 1253.890 1401.100 ;
        RECT 1252.650 1400.900 1253.890 1401.040 ;
        RECT 1252.650 1400.840 1252.970 1400.900 ;
        RECT 1253.570 1400.840 1253.890 1400.900 ;
        RECT 1251.270 1365.680 1251.590 1365.740 ;
        RECT 1253.570 1365.680 1253.890 1365.740 ;
        RECT 1251.270 1365.540 1253.890 1365.680 ;
        RECT 1251.270 1365.480 1251.590 1365.540 ;
        RECT 1253.570 1365.480 1253.890 1365.540 ;
        RECT 1252.190 1304.140 1252.510 1304.200 ;
        RECT 1253.585 1304.140 1253.875 1304.185 ;
        RECT 1252.190 1304.000 1253.875 1304.140 ;
        RECT 1252.190 1303.940 1252.510 1304.000 ;
        RECT 1253.585 1303.955 1253.875 1304.000 ;
        RECT 1253.570 1269.120 1253.890 1269.180 ;
        RECT 1253.375 1268.980 1253.890 1269.120 ;
        RECT 1253.570 1268.920 1253.890 1268.980 ;
        RECT 1253.570 1173.040 1253.890 1173.300 ;
        RECT 1253.660 1172.620 1253.800 1173.040 ;
        RECT 1253.570 1172.360 1253.890 1172.620 ;
        RECT 1252.665 703.700 1252.955 703.745 ;
        RECT 1253.110 703.700 1253.430 703.760 ;
        RECT 1252.665 703.560 1253.430 703.700 ;
        RECT 1252.665 703.515 1252.955 703.560 ;
        RECT 1253.110 703.500 1253.430 703.560 ;
        RECT 1252.650 641.480 1252.970 641.540 ;
        RECT 1252.455 641.340 1252.970 641.480 ;
        RECT 1252.650 641.280 1252.970 641.340 ;
        RECT 1253.110 627.540 1253.430 627.600 ;
        RECT 1253.570 627.540 1253.890 627.600 ;
        RECT 1253.110 627.400 1253.890 627.540 ;
        RECT 1253.110 627.340 1253.430 627.400 ;
        RECT 1253.570 627.340 1253.890 627.400 ;
        RECT 1253.125 558.860 1253.415 558.905 ;
        RECT 1253.570 558.860 1253.890 558.920 ;
        RECT 1253.125 558.720 1253.890 558.860 ;
        RECT 1253.125 558.675 1253.415 558.720 ;
        RECT 1253.570 558.660 1253.890 558.720 ;
        RECT 1253.110 510.920 1253.430 510.980 ;
        RECT 1252.915 510.780 1253.430 510.920 ;
        RECT 1253.110 510.720 1253.430 510.780 ;
        RECT 1253.110 414.020 1253.430 414.080 ;
        RECT 1253.585 414.020 1253.875 414.065 ;
        RECT 1253.110 413.880 1253.875 414.020 ;
        RECT 1253.110 413.820 1253.430 413.880 ;
        RECT 1253.585 413.835 1253.875 413.880 ;
        RECT 1252.190 341.600 1252.510 341.660 ;
        RECT 1253.585 341.600 1253.875 341.645 ;
        RECT 1252.190 341.460 1253.875 341.600 ;
        RECT 1252.190 341.400 1252.510 341.460 ;
        RECT 1253.585 341.415 1253.875 341.460 ;
        RECT 1252.205 96.460 1252.495 96.505 ;
        RECT 1252.650 96.460 1252.970 96.520 ;
        RECT 1252.205 96.320 1252.970 96.460 ;
        RECT 1252.205 96.275 1252.495 96.320 ;
        RECT 1252.650 96.260 1252.970 96.320 ;
        RECT 1252.190 48.520 1252.510 48.580 ;
        RECT 1251.995 48.380 1252.510 48.520 ;
        RECT 1252.190 48.320 1252.510 48.380 ;
        RECT 1001.950 41.380 1002.270 41.440 ;
        RECT 1252.650 41.380 1252.970 41.440 ;
        RECT 1001.950 41.240 1252.970 41.380 ;
        RECT 1001.950 41.180 1002.270 41.240 ;
        RECT 1252.650 41.180 1252.970 41.240 ;
      LAYER via ;
        RECT 1252.680 1666.380 1252.940 1666.640 ;
        RECT 1253.140 1642.240 1253.400 1642.500 ;
        RECT 1252.680 1400.840 1252.940 1401.100 ;
        RECT 1253.600 1400.840 1253.860 1401.100 ;
        RECT 1251.300 1365.480 1251.560 1365.740 ;
        RECT 1253.600 1365.480 1253.860 1365.740 ;
        RECT 1252.220 1303.940 1252.480 1304.200 ;
        RECT 1253.600 1268.920 1253.860 1269.180 ;
        RECT 1253.600 1173.040 1253.860 1173.300 ;
        RECT 1253.600 1172.360 1253.860 1172.620 ;
        RECT 1253.140 703.500 1253.400 703.760 ;
        RECT 1252.680 641.280 1252.940 641.540 ;
        RECT 1253.140 627.340 1253.400 627.600 ;
        RECT 1253.600 627.340 1253.860 627.600 ;
        RECT 1253.600 558.660 1253.860 558.920 ;
        RECT 1253.140 510.720 1253.400 510.980 ;
        RECT 1253.140 413.820 1253.400 414.080 ;
        RECT 1252.220 341.400 1252.480 341.660 ;
        RECT 1252.680 96.260 1252.940 96.520 ;
        RECT 1252.220 48.320 1252.480 48.580 ;
        RECT 1001.980 41.180 1002.240 41.440 ;
        RECT 1252.680 41.180 1252.940 41.440 ;
      LAYER met2 ;
        RECT 1252.580 1700.340 1252.860 1704.000 ;
        RECT 1252.580 1700.000 1252.880 1700.340 ;
        RECT 1252.740 1666.670 1252.880 1700.000 ;
        RECT 1252.680 1666.350 1252.940 1666.670 ;
        RECT 1253.140 1642.210 1253.400 1642.530 ;
        RECT 1253.200 1558.970 1253.340 1642.210 ;
        RECT 1253.200 1558.830 1253.800 1558.970 ;
        RECT 1253.660 1401.130 1253.800 1558.830 ;
        RECT 1252.680 1400.810 1252.940 1401.130 ;
        RECT 1253.600 1400.810 1253.860 1401.130 ;
        RECT 1251.290 1400.275 1251.570 1400.645 ;
        RECT 1252.210 1400.530 1252.490 1400.645 ;
        RECT 1252.740 1400.530 1252.880 1400.810 ;
        RECT 1252.210 1400.390 1252.880 1400.530 ;
        RECT 1252.210 1400.275 1252.490 1400.390 ;
        RECT 1251.360 1365.770 1251.500 1400.275 ;
        RECT 1251.300 1365.450 1251.560 1365.770 ;
        RECT 1253.600 1365.450 1253.860 1365.770 ;
        RECT 1253.660 1305.445 1253.800 1365.450 ;
        RECT 1253.590 1305.075 1253.870 1305.445 ;
        RECT 1252.210 1304.395 1252.490 1304.765 ;
        RECT 1252.280 1304.230 1252.420 1304.395 ;
        RECT 1252.220 1303.910 1252.480 1304.230 ;
        RECT 1253.600 1268.890 1253.860 1269.210 ;
        RECT 1253.660 1173.330 1253.800 1268.890 ;
        RECT 1253.600 1173.010 1253.860 1173.330 ;
        RECT 1253.600 1172.330 1253.860 1172.650 ;
        RECT 1253.660 1125.130 1253.800 1172.330 ;
        RECT 1253.200 1124.990 1253.800 1125.130 ;
        RECT 1253.200 1124.450 1253.340 1124.990 ;
        RECT 1253.200 1124.310 1253.800 1124.450 ;
        RECT 1253.660 1028.570 1253.800 1124.310 ;
        RECT 1253.200 1028.430 1253.800 1028.570 ;
        RECT 1253.200 1027.890 1253.340 1028.430 ;
        RECT 1253.200 1027.750 1253.800 1027.890 ;
        RECT 1253.660 932.010 1253.800 1027.750 ;
        RECT 1253.200 931.870 1253.800 932.010 ;
        RECT 1253.200 931.330 1253.340 931.870 ;
        RECT 1253.200 931.190 1253.800 931.330 ;
        RECT 1253.660 835.450 1253.800 931.190 ;
        RECT 1253.200 835.310 1253.800 835.450 ;
        RECT 1253.200 834.770 1253.340 835.310 ;
        RECT 1253.200 834.630 1253.800 834.770 ;
        RECT 1253.660 711.805 1253.800 834.630 ;
        RECT 1253.590 711.435 1253.870 711.805 ;
        RECT 1253.130 710.755 1253.410 711.125 ;
        RECT 1253.200 703.790 1253.340 710.755 ;
        RECT 1253.140 703.470 1253.400 703.790 ;
        RECT 1252.680 641.250 1252.940 641.570 ;
        RECT 1252.740 628.050 1252.880 641.250 ;
        RECT 1252.740 627.910 1253.340 628.050 ;
        RECT 1253.200 627.630 1253.340 627.910 ;
        RECT 1253.140 627.310 1253.400 627.630 ;
        RECT 1253.600 627.310 1253.860 627.630 ;
        RECT 1253.660 558.950 1253.800 627.310 ;
        RECT 1253.600 558.630 1253.860 558.950 ;
        RECT 1253.140 510.690 1253.400 511.010 ;
        RECT 1253.200 414.110 1253.340 510.690 ;
        RECT 1253.140 413.790 1253.400 414.110 ;
        RECT 1252.220 341.370 1252.480 341.690 ;
        RECT 1252.280 290.090 1252.420 341.370 ;
        RECT 1252.280 289.950 1252.880 290.090 ;
        RECT 1252.740 241.810 1252.880 289.950 ;
        RECT 1252.280 241.670 1252.880 241.810 ;
        RECT 1252.280 220.845 1252.420 241.670 ;
        RECT 1252.210 220.475 1252.490 220.845 ;
        RECT 1253.590 220.475 1253.870 220.845 ;
        RECT 1253.660 96.970 1253.800 220.475 ;
        RECT 1252.740 96.830 1253.800 96.970 ;
        RECT 1252.740 96.550 1252.880 96.830 ;
        RECT 1252.680 96.230 1252.940 96.550 ;
        RECT 1252.220 48.290 1252.480 48.610 ;
        RECT 1252.280 48.010 1252.420 48.290 ;
        RECT 1252.280 47.870 1252.880 48.010 ;
        RECT 1252.740 41.470 1252.880 47.870 ;
        RECT 1001.980 41.150 1002.240 41.470 ;
        RECT 1252.680 41.150 1252.940 41.470 ;
        RECT 1002.040 2.400 1002.180 41.150 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
      LAYER via2 ;
        RECT 1251.290 1400.320 1251.570 1400.600 ;
        RECT 1252.210 1400.320 1252.490 1400.600 ;
        RECT 1253.590 1305.120 1253.870 1305.400 ;
        RECT 1252.210 1304.440 1252.490 1304.720 ;
        RECT 1253.590 711.480 1253.870 711.760 ;
        RECT 1253.130 710.800 1253.410 711.080 ;
        RECT 1252.210 220.520 1252.490 220.800 ;
        RECT 1253.590 220.520 1253.870 220.800 ;
      LAYER met3 ;
        RECT 1251.265 1400.610 1251.595 1400.625 ;
        RECT 1252.185 1400.610 1252.515 1400.625 ;
        RECT 1251.265 1400.310 1252.515 1400.610 ;
        RECT 1251.265 1400.295 1251.595 1400.310 ;
        RECT 1252.185 1400.295 1252.515 1400.310 ;
        RECT 1253.565 1305.410 1253.895 1305.425 ;
        RECT 1251.510 1305.110 1253.895 1305.410 ;
        RECT 1251.510 1304.730 1251.810 1305.110 ;
        RECT 1253.565 1305.095 1253.895 1305.110 ;
        RECT 1252.185 1304.730 1252.515 1304.745 ;
        RECT 1251.510 1304.430 1252.515 1304.730 ;
        RECT 1252.185 1304.415 1252.515 1304.430 ;
        RECT 1253.565 711.770 1253.895 711.785 ;
        RECT 1252.430 711.470 1253.895 711.770 ;
        RECT 1252.430 711.090 1252.730 711.470 ;
        RECT 1253.565 711.455 1253.895 711.470 ;
        RECT 1253.105 711.090 1253.435 711.105 ;
        RECT 1252.430 710.790 1253.435 711.090 ;
        RECT 1253.105 710.775 1253.435 710.790 ;
        RECT 1252.185 220.810 1252.515 220.825 ;
        RECT 1253.565 220.810 1253.895 220.825 ;
        RECT 1252.185 220.510 1253.895 220.810 ;
        RECT 1252.185 220.495 1252.515 220.510 ;
        RECT 1253.565 220.495 1253.895 220.510 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1254.565 362.185 1254.735 386.155 ;
      LAYER mcon ;
        RECT 1254.565 385.985 1254.735 386.155 ;
      LAYER met1 ;
        RECT 1254.490 386.140 1254.810 386.200 ;
        RECT 1254.295 386.000 1254.810 386.140 ;
        RECT 1254.490 385.940 1254.810 386.000 ;
        RECT 1254.490 362.340 1254.810 362.400 ;
        RECT 1254.295 362.200 1254.810 362.340 ;
        RECT 1254.490 362.140 1254.810 362.200 ;
        RECT 1019.430 37.640 1019.750 37.700 ;
        RECT 1254.490 37.640 1254.810 37.700 ;
        RECT 1019.430 37.500 1254.810 37.640 ;
        RECT 1019.430 37.440 1019.750 37.500 ;
        RECT 1254.490 37.440 1254.810 37.500 ;
      LAYER via ;
        RECT 1254.520 385.940 1254.780 386.200 ;
        RECT 1254.520 362.140 1254.780 362.400 ;
        RECT 1019.460 37.440 1019.720 37.700 ;
        RECT 1254.520 37.440 1254.780 37.700 ;
      LAYER met2 ;
        RECT 1254.420 1700.340 1254.700 1704.000 ;
        RECT 1254.420 1700.000 1254.720 1700.340 ;
        RECT 1254.580 386.230 1254.720 1700.000 ;
        RECT 1254.520 385.910 1254.780 386.230 ;
        RECT 1254.520 362.110 1254.780 362.430 ;
        RECT 1254.580 37.730 1254.720 362.110 ;
        RECT 1019.460 37.410 1019.720 37.730 ;
        RECT 1254.520 37.410 1254.780 37.730 ;
        RECT 1019.520 2.400 1019.660 37.410 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1242.530 1684.940 1242.850 1685.000 ;
        RECT 1256.330 1684.940 1256.650 1685.000 ;
        RECT 1242.530 1684.800 1256.650 1684.940 ;
        RECT 1242.530 1684.740 1242.850 1684.800 ;
        RECT 1256.330 1684.740 1256.650 1684.800 ;
        RECT 1041.510 1654.000 1041.830 1654.060 ;
        RECT 1242.070 1654.000 1242.390 1654.060 ;
        RECT 1041.510 1653.860 1242.390 1654.000 ;
        RECT 1041.510 1653.800 1041.830 1653.860 ;
        RECT 1242.070 1653.800 1242.390 1653.860 ;
        RECT 1037.370 2.960 1037.690 3.020 ;
        RECT 1041.510 2.960 1041.830 3.020 ;
        RECT 1037.370 2.820 1041.830 2.960 ;
        RECT 1037.370 2.760 1037.690 2.820 ;
        RECT 1041.510 2.760 1041.830 2.820 ;
      LAYER via ;
        RECT 1242.560 1684.740 1242.820 1685.000 ;
        RECT 1256.360 1684.740 1256.620 1685.000 ;
        RECT 1041.540 1653.800 1041.800 1654.060 ;
        RECT 1242.100 1653.800 1242.360 1654.060 ;
        RECT 1037.400 2.760 1037.660 3.020 ;
        RECT 1041.540 2.760 1041.800 3.020 ;
      LAYER met2 ;
        RECT 1256.260 1700.340 1256.540 1704.000 ;
        RECT 1256.260 1700.000 1256.560 1700.340 ;
        RECT 1256.420 1685.030 1256.560 1700.000 ;
        RECT 1242.560 1684.710 1242.820 1685.030 ;
        RECT 1256.360 1684.710 1256.620 1685.030 ;
        RECT 1242.620 1677.970 1242.760 1684.710 ;
        RECT 1242.160 1677.830 1242.760 1677.970 ;
        RECT 1242.160 1654.090 1242.300 1677.830 ;
        RECT 1041.540 1653.770 1041.800 1654.090 ;
        RECT 1242.100 1653.770 1242.360 1654.090 ;
        RECT 1041.600 3.050 1041.740 1653.770 ;
        RECT 1037.400 2.730 1037.660 3.050 ;
        RECT 1041.540 2.730 1041.800 3.050 ;
        RECT 1037.460 2.400 1037.600 2.730 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1258.170 1676.240 1258.490 1676.500 ;
        RECT 1258.260 1675.420 1258.400 1676.240 ;
        RECT 1258.630 1675.420 1258.950 1675.480 ;
        RECT 1258.260 1675.280 1258.950 1675.420 ;
        RECT 1258.630 1675.220 1258.950 1675.280 ;
        RECT 1054.850 1597.900 1055.170 1597.960 ;
        RECT 1258.630 1597.900 1258.950 1597.960 ;
        RECT 1054.850 1597.760 1258.950 1597.900 ;
        RECT 1054.850 1597.700 1055.170 1597.760 ;
        RECT 1258.630 1597.700 1258.950 1597.760 ;
      LAYER via ;
        RECT 1258.200 1676.240 1258.460 1676.500 ;
        RECT 1258.660 1675.220 1258.920 1675.480 ;
        RECT 1054.880 1597.700 1055.140 1597.960 ;
        RECT 1258.660 1597.700 1258.920 1597.960 ;
      LAYER met2 ;
        RECT 1258.100 1700.340 1258.380 1704.000 ;
        RECT 1258.100 1700.000 1258.400 1700.340 ;
        RECT 1258.260 1676.530 1258.400 1700.000 ;
        RECT 1258.200 1676.210 1258.460 1676.530 ;
        RECT 1258.660 1675.190 1258.920 1675.510 ;
        RECT 1258.720 1597.990 1258.860 1675.190 ;
        RECT 1054.880 1597.670 1055.140 1597.990 ;
        RECT 1258.660 1597.670 1258.920 1597.990 ;
        RECT 1054.940 17.410 1055.080 1597.670 ;
        RECT 1054.940 17.270 1055.540 17.410 ;
        RECT 1055.400 2.400 1055.540 17.270 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1076.010 1640.060 1076.330 1640.120 ;
        RECT 1258.170 1640.060 1258.490 1640.120 ;
        RECT 1076.010 1639.920 1258.490 1640.060 ;
        RECT 1076.010 1639.860 1076.330 1639.920 ;
        RECT 1258.170 1639.860 1258.490 1639.920 ;
      LAYER via ;
        RECT 1076.040 1639.860 1076.300 1640.120 ;
        RECT 1258.200 1639.860 1258.460 1640.120 ;
      LAYER met2 ;
        RECT 1259.940 1700.340 1260.220 1704.000 ;
        RECT 1259.940 1700.000 1260.240 1700.340 ;
        RECT 1260.100 1675.930 1260.240 1700.000 ;
        RECT 1258.260 1675.790 1260.240 1675.930 ;
        RECT 1258.260 1640.150 1258.400 1675.790 ;
        RECT 1076.040 1639.830 1076.300 1640.150 ;
        RECT 1258.200 1639.830 1258.460 1640.150 ;
        RECT 1076.100 18.090 1076.240 1639.830 ;
        RECT 1073.340 17.950 1076.240 18.090 ;
        RECT 1073.340 2.400 1073.480 17.950 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1261.005 1248.905 1261.175 1256.555 ;
        RECT 1261.005 993.565 1261.175 1041.675 ;
        RECT 1260.545 883.405 1260.715 931.515 ;
        RECT 1261.005 841.585 1261.175 869.975 ;
      LAYER mcon ;
        RECT 1261.005 1256.385 1261.175 1256.555 ;
        RECT 1261.005 1041.505 1261.175 1041.675 ;
        RECT 1260.545 931.345 1260.715 931.515 ;
        RECT 1261.005 869.805 1261.175 869.975 ;
      LAYER met1 ;
        RECT 1259.550 1669.980 1259.870 1670.040 ;
        RECT 1261.850 1669.980 1262.170 1670.040 ;
        RECT 1259.550 1669.840 1262.170 1669.980 ;
        RECT 1259.550 1669.780 1259.870 1669.840 ;
        RECT 1261.850 1669.780 1262.170 1669.840 ;
        RECT 1259.550 1631.900 1259.870 1631.960 ;
        RECT 1260.470 1631.900 1260.790 1631.960 ;
        RECT 1259.550 1631.760 1260.790 1631.900 ;
        RECT 1259.550 1631.700 1259.870 1631.760 ;
        RECT 1260.470 1631.700 1260.790 1631.760 ;
        RECT 1260.930 1483.320 1261.250 1483.380 ;
        RECT 1261.390 1483.320 1261.710 1483.380 ;
        RECT 1260.930 1483.180 1261.710 1483.320 ;
        RECT 1260.930 1483.120 1261.250 1483.180 ;
        RECT 1261.390 1483.120 1261.710 1483.180 ;
        RECT 1260.945 1256.540 1261.235 1256.585 ;
        RECT 1261.390 1256.540 1261.710 1256.600 ;
        RECT 1260.945 1256.400 1261.710 1256.540 ;
        RECT 1260.945 1256.355 1261.235 1256.400 ;
        RECT 1261.390 1256.340 1261.710 1256.400 ;
        RECT 1260.930 1249.060 1261.250 1249.120 ;
        RECT 1260.735 1248.920 1261.250 1249.060 ;
        RECT 1260.930 1248.860 1261.250 1248.920 ;
        RECT 1260.470 1221.180 1260.790 1221.240 ;
        RECT 1261.390 1221.180 1261.710 1221.240 ;
        RECT 1260.470 1221.040 1261.710 1221.180 ;
        RECT 1260.470 1220.980 1260.790 1221.040 ;
        RECT 1261.390 1220.980 1261.710 1221.040 ;
        RECT 1260.930 1041.660 1261.250 1041.720 ;
        RECT 1260.735 1041.520 1261.250 1041.660 ;
        RECT 1260.930 1041.460 1261.250 1041.520 ;
        RECT 1260.945 993.720 1261.235 993.765 ;
        RECT 1261.390 993.720 1261.710 993.780 ;
        RECT 1260.945 993.580 1261.710 993.720 ;
        RECT 1260.945 993.535 1261.235 993.580 ;
        RECT 1261.390 993.520 1261.710 993.580 ;
        RECT 1260.470 945.440 1260.790 945.500 ;
        RECT 1261.390 945.440 1261.710 945.500 ;
        RECT 1260.470 945.300 1261.710 945.440 ;
        RECT 1260.470 945.240 1260.790 945.300 ;
        RECT 1261.390 945.240 1261.710 945.300 ;
        RECT 1260.470 931.500 1260.790 931.560 ;
        RECT 1260.275 931.360 1260.790 931.500 ;
        RECT 1260.470 931.300 1260.790 931.360 ;
        RECT 1260.485 883.560 1260.775 883.605 ;
        RECT 1260.930 883.560 1261.250 883.620 ;
        RECT 1260.485 883.420 1261.250 883.560 ;
        RECT 1260.485 883.375 1260.775 883.420 ;
        RECT 1260.930 883.360 1261.250 883.420 ;
        RECT 1260.930 869.960 1261.250 870.020 ;
        RECT 1260.735 869.820 1261.250 869.960 ;
        RECT 1260.930 869.760 1261.250 869.820 ;
        RECT 1260.930 841.740 1261.250 841.800 ;
        RECT 1260.735 841.600 1261.250 841.740 ;
        RECT 1260.930 841.540 1261.250 841.600 ;
        RECT 1096.250 824.400 1096.570 824.460 ;
        RECT 1260.930 824.400 1261.250 824.460 ;
        RECT 1096.250 824.260 1261.250 824.400 ;
        RECT 1096.250 824.200 1096.570 824.260 ;
        RECT 1260.930 824.200 1261.250 824.260 ;
      LAYER via ;
        RECT 1259.580 1669.780 1259.840 1670.040 ;
        RECT 1261.880 1669.780 1262.140 1670.040 ;
        RECT 1259.580 1631.700 1259.840 1631.960 ;
        RECT 1260.500 1631.700 1260.760 1631.960 ;
        RECT 1260.960 1483.120 1261.220 1483.380 ;
        RECT 1261.420 1483.120 1261.680 1483.380 ;
        RECT 1261.420 1256.340 1261.680 1256.600 ;
        RECT 1260.960 1248.860 1261.220 1249.120 ;
        RECT 1260.500 1220.980 1260.760 1221.240 ;
        RECT 1261.420 1220.980 1261.680 1221.240 ;
        RECT 1260.960 1041.460 1261.220 1041.720 ;
        RECT 1261.420 993.520 1261.680 993.780 ;
        RECT 1260.500 945.240 1260.760 945.500 ;
        RECT 1261.420 945.240 1261.680 945.500 ;
        RECT 1260.500 931.300 1260.760 931.560 ;
        RECT 1260.960 883.360 1261.220 883.620 ;
        RECT 1260.960 869.760 1261.220 870.020 ;
        RECT 1260.960 841.540 1261.220 841.800 ;
        RECT 1096.280 824.200 1096.540 824.460 ;
        RECT 1260.960 824.200 1261.220 824.460 ;
      LAYER met2 ;
        RECT 1261.780 1700.340 1262.060 1704.000 ;
        RECT 1261.780 1700.000 1262.080 1700.340 ;
        RECT 1261.940 1670.070 1262.080 1700.000 ;
        RECT 1259.580 1669.750 1259.840 1670.070 ;
        RECT 1261.880 1669.750 1262.140 1670.070 ;
        RECT 1259.640 1631.990 1259.780 1669.750 ;
        RECT 1259.580 1631.670 1259.840 1631.990 ;
        RECT 1260.500 1631.670 1260.760 1631.990 ;
        RECT 1260.560 1558.970 1260.700 1631.670 ;
        RECT 1260.560 1558.830 1261.160 1558.970 ;
        RECT 1261.020 1483.410 1261.160 1558.830 ;
        RECT 1260.960 1483.090 1261.220 1483.410 ;
        RECT 1261.420 1483.090 1261.680 1483.410 ;
        RECT 1261.480 1256.630 1261.620 1483.090 ;
        RECT 1261.420 1256.310 1261.680 1256.630 ;
        RECT 1260.960 1248.830 1261.220 1249.150 ;
        RECT 1261.020 1221.690 1261.160 1248.830 ;
        RECT 1260.560 1221.550 1261.160 1221.690 ;
        RECT 1260.560 1221.270 1260.700 1221.550 ;
        RECT 1260.500 1220.950 1260.760 1221.270 ;
        RECT 1261.420 1220.950 1261.680 1221.270 ;
        RECT 1261.480 1145.530 1261.620 1220.950 ;
        RECT 1261.020 1145.390 1261.620 1145.530 ;
        RECT 1261.020 1041.750 1261.160 1145.390 ;
        RECT 1260.960 1041.430 1261.220 1041.750 ;
        RECT 1261.420 993.490 1261.680 993.810 ;
        RECT 1261.480 945.530 1261.620 993.490 ;
        RECT 1260.500 945.210 1260.760 945.530 ;
        RECT 1261.420 945.210 1261.680 945.530 ;
        RECT 1260.560 931.590 1260.700 945.210 ;
        RECT 1260.500 931.270 1260.760 931.590 ;
        RECT 1260.960 883.330 1261.220 883.650 ;
        RECT 1261.020 870.050 1261.160 883.330 ;
        RECT 1260.960 869.730 1261.220 870.050 ;
        RECT 1260.960 841.510 1261.220 841.830 ;
        RECT 1261.020 824.490 1261.160 841.510 ;
        RECT 1096.280 824.170 1096.540 824.490 ;
        RECT 1260.960 824.170 1261.220 824.490 ;
        RECT 1096.340 18.090 1096.480 824.170 ;
        RECT 1090.820 17.950 1096.480 18.090 ;
        RECT 1090.820 2.400 1090.960 17.950 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1110.510 1633.260 1110.830 1633.320 ;
        RECT 1263.690 1633.260 1264.010 1633.320 ;
        RECT 1110.510 1633.120 1264.010 1633.260 ;
        RECT 1110.510 1633.060 1110.830 1633.120 ;
        RECT 1263.690 1633.060 1264.010 1633.120 ;
      LAYER via ;
        RECT 1110.540 1633.060 1110.800 1633.320 ;
        RECT 1263.720 1633.060 1263.980 1633.320 ;
      LAYER met2 ;
        RECT 1263.620 1700.340 1263.900 1704.000 ;
        RECT 1263.620 1700.000 1263.920 1700.340 ;
        RECT 1263.780 1633.350 1263.920 1700.000 ;
        RECT 1110.540 1633.030 1110.800 1633.350 ;
        RECT 1263.720 1633.030 1263.980 1633.350 ;
        RECT 1110.600 16.730 1110.740 1633.030 ;
        RECT 1108.760 16.590 1110.740 16.730 ;
        RECT 1108.760 2.400 1108.900 16.590 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1131.210 1612.180 1131.530 1612.240 ;
        RECT 1265.530 1612.180 1265.850 1612.240 ;
        RECT 1131.210 1612.040 1265.850 1612.180 ;
        RECT 1131.210 1611.980 1131.530 1612.040 ;
        RECT 1265.530 1611.980 1265.850 1612.040 ;
        RECT 1126.610 19.280 1126.930 19.340 ;
        RECT 1131.210 19.280 1131.530 19.340 ;
        RECT 1126.610 19.140 1131.530 19.280 ;
        RECT 1126.610 19.080 1126.930 19.140 ;
        RECT 1131.210 19.080 1131.530 19.140 ;
      LAYER via ;
        RECT 1131.240 1611.980 1131.500 1612.240 ;
        RECT 1265.560 1611.980 1265.820 1612.240 ;
        RECT 1126.640 19.080 1126.900 19.340 ;
        RECT 1131.240 19.080 1131.500 19.340 ;
      LAYER met2 ;
        RECT 1265.460 1700.340 1265.740 1704.000 ;
        RECT 1265.460 1700.000 1265.760 1700.340 ;
        RECT 1265.620 1612.270 1265.760 1700.000 ;
        RECT 1131.240 1611.950 1131.500 1612.270 ;
        RECT 1265.560 1611.950 1265.820 1612.270 ;
        RECT 1131.300 19.370 1131.440 1611.950 ;
        RECT 1126.640 19.050 1126.900 19.370 ;
        RECT 1131.240 19.050 1131.500 19.370 ;
        RECT 1126.700 2.400 1126.840 19.050 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1260.010 1642.440 1260.330 1642.500 ;
        RECT 1267.370 1642.440 1267.690 1642.500 ;
        RECT 1260.010 1642.300 1267.690 1642.440 ;
        RECT 1260.010 1642.240 1260.330 1642.300 ;
        RECT 1267.370 1642.240 1267.690 1642.300 ;
        RECT 1144.550 58.720 1144.870 58.780 ;
        RECT 1260.010 58.720 1260.330 58.780 ;
        RECT 1144.550 58.580 1260.330 58.720 ;
        RECT 1144.550 58.520 1144.870 58.580 ;
        RECT 1260.010 58.520 1260.330 58.580 ;
      LAYER via ;
        RECT 1260.040 1642.240 1260.300 1642.500 ;
        RECT 1267.400 1642.240 1267.660 1642.500 ;
        RECT 1144.580 58.520 1144.840 58.780 ;
        RECT 1260.040 58.520 1260.300 58.780 ;
      LAYER met2 ;
        RECT 1267.300 1700.340 1267.580 1704.000 ;
        RECT 1267.300 1700.000 1267.600 1700.340 ;
        RECT 1267.460 1642.530 1267.600 1700.000 ;
        RECT 1260.040 1642.210 1260.300 1642.530 ;
        RECT 1267.400 1642.210 1267.660 1642.530 ;
        RECT 1260.100 58.810 1260.240 1642.210 ;
        RECT 1144.580 58.490 1144.840 58.810 ;
        RECT 1260.040 58.490 1260.300 58.810 ;
        RECT 1144.640 2.400 1144.780 58.490 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1264.610 1678.140 1264.930 1678.200 ;
        RECT 1269.210 1678.140 1269.530 1678.200 ;
        RECT 1264.610 1678.000 1269.530 1678.140 ;
        RECT 1264.610 1677.940 1264.930 1678.000 ;
        RECT 1269.210 1677.940 1269.530 1678.000 ;
        RECT 1162.490 51.920 1162.810 51.980 ;
        RECT 1264.610 51.920 1264.930 51.980 ;
        RECT 1162.490 51.780 1264.930 51.920 ;
        RECT 1162.490 51.720 1162.810 51.780 ;
        RECT 1264.610 51.720 1264.930 51.780 ;
      LAYER via ;
        RECT 1264.640 1677.940 1264.900 1678.200 ;
        RECT 1269.240 1677.940 1269.500 1678.200 ;
        RECT 1162.520 51.720 1162.780 51.980 ;
        RECT 1264.640 51.720 1264.900 51.980 ;
      LAYER met2 ;
        RECT 1269.140 1700.340 1269.420 1704.000 ;
        RECT 1269.140 1700.000 1269.440 1700.340 ;
        RECT 1269.300 1678.230 1269.440 1700.000 ;
        RECT 1264.640 1677.910 1264.900 1678.230 ;
        RECT 1269.240 1677.910 1269.500 1678.230 ;
        RECT 1264.700 52.010 1264.840 1677.910 ;
        RECT 1162.520 51.690 1162.780 52.010 ;
        RECT 1264.640 51.690 1264.900 52.010 ;
        RECT 1162.580 2.400 1162.720 51.690 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 682.710 1591.100 683.030 1591.160 ;
        RECT 1219.530 1591.100 1219.850 1591.160 ;
        RECT 682.710 1590.960 1219.850 1591.100 ;
        RECT 682.710 1590.900 683.030 1590.960 ;
        RECT 1219.530 1590.900 1219.850 1590.960 ;
      LAYER via ;
        RECT 682.740 1590.900 683.000 1591.160 ;
        RECT 1219.560 1590.900 1219.820 1591.160 ;
      LAYER met2 ;
        RECT 1219.460 1700.340 1219.740 1704.000 ;
        RECT 1219.460 1700.000 1219.760 1700.340 ;
        RECT 1219.620 1591.190 1219.760 1700.000 ;
        RECT 682.740 1590.870 683.000 1591.190 ;
        RECT 1219.560 1590.870 1219.820 1591.190 ;
        RECT 682.800 24.210 682.940 1590.870 ;
        RECT 680.500 24.070 682.940 24.210 ;
        RECT 680.500 2.400 680.640 24.070 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1265.990 1689.700 1266.310 1689.760 ;
        RECT 1271.050 1689.700 1271.370 1689.760 ;
        RECT 1265.990 1689.560 1271.370 1689.700 ;
        RECT 1265.990 1689.500 1266.310 1689.560 ;
        RECT 1271.050 1689.500 1271.370 1689.560 ;
        RECT 1179.970 52.260 1180.290 52.320 ;
        RECT 1265.990 52.260 1266.310 52.320 ;
        RECT 1179.970 52.120 1266.310 52.260 ;
        RECT 1179.970 52.060 1180.290 52.120 ;
        RECT 1265.990 52.060 1266.310 52.120 ;
      LAYER via ;
        RECT 1266.020 1689.500 1266.280 1689.760 ;
        RECT 1271.080 1689.500 1271.340 1689.760 ;
        RECT 1180.000 52.060 1180.260 52.320 ;
        RECT 1266.020 52.060 1266.280 52.320 ;
      LAYER met2 ;
        RECT 1270.980 1700.340 1271.260 1704.000 ;
        RECT 1270.980 1700.000 1271.280 1700.340 ;
        RECT 1271.140 1689.790 1271.280 1700.000 ;
        RECT 1266.020 1689.470 1266.280 1689.790 ;
        RECT 1271.080 1689.470 1271.340 1689.790 ;
        RECT 1266.080 52.350 1266.220 1689.470 ;
        RECT 1180.000 52.030 1180.260 52.350 ;
        RECT 1266.020 52.030 1266.280 52.350 ;
        RECT 1180.060 2.400 1180.200 52.030 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1200.285 1676.965 1200.455 1685.635 ;
      LAYER mcon ;
        RECT 1200.285 1685.465 1200.455 1685.635 ;
      LAYER met1 ;
        RECT 1200.225 1685.620 1200.515 1685.665 ;
        RECT 1272.890 1685.620 1273.210 1685.680 ;
        RECT 1200.225 1685.480 1273.210 1685.620 ;
        RECT 1200.225 1685.435 1200.515 1685.480 ;
        RECT 1272.890 1685.420 1273.210 1685.480 ;
        RECT 1200.210 1677.120 1200.530 1677.180 ;
        RECT 1200.015 1676.980 1200.530 1677.120 ;
        RECT 1200.210 1676.920 1200.530 1676.980 ;
        RECT 1197.910 20.640 1198.230 20.700 ;
        RECT 1200.210 20.640 1200.530 20.700 ;
        RECT 1197.910 20.500 1200.530 20.640 ;
        RECT 1197.910 20.440 1198.230 20.500 ;
        RECT 1200.210 20.440 1200.530 20.500 ;
      LAYER via ;
        RECT 1272.920 1685.420 1273.180 1685.680 ;
        RECT 1200.240 1676.920 1200.500 1677.180 ;
        RECT 1197.940 20.440 1198.200 20.700 ;
        RECT 1200.240 20.440 1200.500 20.700 ;
      LAYER met2 ;
        RECT 1272.820 1700.340 1273.100 1704.000 ;
        RECT 1272.820 1700.000 1273.120 1700.340 ;
        RECT 1272.980 1685.710 1273.120 1700.000 ;
        RECT 1272.920 1685.390 1273.180 1685.710 ;
        RECT 1200.240 1676.890 1200.500 1677.210 ;
        RECT 1200.300 20.730 1200.440 1676.890 ;
        RECT 1197.940 20.410 1198.200 20.730 ;
        RECT 1200.240 20.410 1200.500 20.730 ;
        RECT 1198.000 2.400 1198.140 20.410 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1274.345 1580.405 1274.515 1669.655 ;
        RECT 1274.345 1428.425 1274.515 1476.535 ;
        RECT 1274.345 1248.905 1274.515 1256.215 ;
        RECT 1273.885 897.005 1274.055 945.115 ;
        RECT 1274.345 793.645 1274.515 841.755 ;
        RECT 1275.265 565.845 1275.435 613.955 ;
        RECT 1274.345 476.085 1274.515 524.195 ;
        RECT 1274.805 255.425 1274.975 303.195 ;
      LAYER mcon ;
        RECT 1274.345 1669.485 1274.515 1669.655 ;
        RECT 1274.345 1476.365 1274.515 1476.535 ;
        RECT 1274.345 1256.045 1274.515 1256.215 ;
        RECT 1273.885 944.945 1274.055 945.115 ;
        RECT 1274.345 841.585 1274.515 841.755 ;
        RECT 1275.265 613.785 1275.435 613.955 ;
        RECT 1274.345 524.025 1274.515 524.195 ;
        RECT 1274.805 303.025 1274.975 303.195 ;
      LAYER met1 ;
        RECT 1274.285 1669.640 1274.575 1669.685 ;
        RECT 1274.730 1669.640 1275.050 1669.700 ;
        RECT 1274.285 1669.500 1275.050 1669.640 ;
        RECT 1274.285 1669.455 1274.575 1669.500 ;
        RECT 1274.730 1669.440 1275.050 1669.500 ;
        RECT 1274.270 1580.560 1274.590 1580.620 ;
        RECT 1274.075 1580.420 1274.590 1580.560 ;
        RECT 1274.270 1580.360 1274.590 1580.420 ;
        RECT 1273.810 1524.800 1274.130 1524.860 ;
        RECT 1275.190 1524.800 1275.510 1524.860 ;
        RECT 1273.810 1524.660 1275.510 1524.800 ;
        RECT 1273.810 1524.600 1274.130 1524.660 ;
        RECT 1275.190 1524.600 1275.510 1524.660 ;
        RECT 1274.270 1476.520 1274.590 1476.580 ;
        RECT 1274.075 1476.380 1274.590 1476.520 ;
        RECT 1274.270 1476.320 1274.590 1476.380 ;
        RECT 1274.270 1428.580 1274.590 1428.640 ;
        RECT 1274.075 1428.440 1274.590 1428.580 ;
        RECT 1274.270 1428.380 1274.590 1428.440 ;
        RECT 1274.270 1256.200 1274.590 1256.260 ;
        RECT 1274.075 1256.060 1274.590 1256.200 ;
        RECT 1274.270 1256.000 1274.590 1256.060 ;
        RECT 1274.270 1249.060 1274.590 1249.120 ;
        RECT 1274.075 1248.920 1274.590 1249.060 ;
        RECT 1274.270 1248.860 1274.590 1248.920 ;
        RECT 1273.810 1110.820 1274.130 1111.080 ;
        RECT 1273.900 1110.680 1274.040 1110.820 ;
        RECT 1274.270 1110.680 1274.590 1110.740 ;
        RECT 1273.900 1110.540 1274.590 1110.680 ;
        RECT 1274.270 1110.480 1274.590 1110.540 ;
        RECT 1274.270 1014.460 1274.590 1014.520 ;
        RECT 1274.730 1014.460 1275.050 1014.520 ;
        RECT 1274.270 1014.320 1275.050 1014.460 ;
        RECT 1274.270 1014.260 1274.590 1014.320 ;
        RECT 1274.730 1014.260 1275.050 1014.320 ;
        RECT 1273.810 945.100 1274.130 945.160 ;
        RECT 1273.615 944.960 1274.130 945.100 ;
        RECT 1273.810 944.900 1274.130 944.960 ;
        RECT 1273.825 897.160 1274.115 897.205 ;
        RECT 1274.730 897.160 1275.050 897.220 ;
        RECT 1273.825 897.020 1275.050 897.160 ;
        RECT 1273.825 896.975 1274.115 897.020 ;
        RECT 1274.730 896.960 1275.050 897.020 ;
        RECT 1274.285 841.740 1274.575 841.785 ;
        RECT 1274.730 841.740 1275.050 841.800 ;
        RECT 1274.285 841.600 1275.050 841.740 ;
        RECT 1274.285 841.555 1274.575 841.600 ;
        RECT 1274.730 841.540 1275.050 841.600 ;
        RECT 1274.270 793.800 1274.590 793.860 ;
        RECT 1274.075 793.660 1274.590 793.800 ;
        RECT 1274.270 793.600 1274.590 793.660 ;
        RECT 1274.270 752.320 1274.590 752.380 ;
        RECT 1275.190 752.320 1275.510 752.380 ;
        RECT 1274.270 752.180 1275.510 752.320 ;
        RECT 1274.270 752.120 1274.590 752.180 ;
        RECT 1275.190 752.120 1275.510 752.180 ;
        RECT 1274.730 703.700 1275.050 703.760 ;
        RECT 1275.190 703.700 1275.510 703.760 ;
        RECT 1274.730 703.560 1275.510 703.700 ;
        RECT 1274.730 703.500 1275.050 703.560 ;
        RECT 1275.190 703.500 1275.510 703.560 ;
        RECT 1274.730 628.220 1275.050 628.280 ;
        RECT 1274.360 628.080 1275.050 628.220 ;
        RECT 1274.360 627.940 1274.500 628.080 ;
        RECT 1274.730 628.020 1275.050 628.080 ;
        RECT 1274.270 627.680 1274.590 627.940 ;
        RECT 1274.270 620.740 1274.590 620.800 ;
        RECT 1275.650 620.740 1275.970 620.800 ;
        RECT 1274.270 620.600 1275.970 620.740 ;
        RECT 1274.270 620.540 1274.590 620.600 ;
        RECT 1275.650 620.540 1275.970 620.600 ;
        RECT 1275.205 613.940 1275.495 613.985 ;
        RECT 1275.650 613.940 1275.970 614.000 ;
        RECT 1275.205 613.800 1275.970 613.940 ;
        RECT 1275.205 613.755 1275.495 613.800 ;
        RECT 1275.650 613.740 1275.970 613.800 ;
        RECT 1275.190 566.000 1275.510 566.060 ;
        RECT 1274.995 565.860 1275.510 566.000 ;
        RECT 1275.190 565.800 1275.510 565.860 ;
        RECT 1274.270 524.180 1274.590 524.240 ;
        RECT 1274.075 524.040 1274.590 524.180 ;
        RECT 1274.270 523.980 1274.590 524.040 ;
        RECT 1274.285 476.240 1274.575 476.285 ;
        RECT 1275.190 476.240 1275.510 476.300 ;
        RECT 1274.285 476.100 1275.510 476.240 ;
        RECT 1274.285 476.055 1274.575 476.100 ;
        RECT 1275.190 476.040 1275.510 476.100 ;
        RECT 1273.810 407.220 1274.130 407.280 ;
        RECT 1274.730 407.220 1275.050 407.280 ;
        RECT 1273.810 407.080 1275.050 407.220 ;
        RECT 1273.810 407.020 1274.130 407.080 ;
        RECT 1274.730 407.020 1275.050 407.080 ;
        RECT 1274.270 303.180 1274.590 303.240 ;
        RECT 1274.745 303.180 1275.035 303.225 ;
        RECT 1274.270 303.040 1275.035 303.180 ;
        RECT 1274.270 302.980 1274.590 303.040 ;
        RECT 1274.745 302.995 1275.035 303.040 ;
        RECT 1274.745 255.580 1275.035 255.625 ;
        RECT 1275.190 255.580 1275.510 255.640 ;
        RECT 1274.745 255.440 1275.510 255.580 ;
        RECT 1274.745 255.395 1275.035 255.440 ;
        RECT 1275.190 255.380 1275.510 255.440 ;
        RECT 1273.810 214.100 1274.130 214.160 ;
        RECT 1275.190 214.100 1275.510 214.160 ;
        RECT 1273.810 213.960 1275.510 214.100 ;
        RECT 1273.810 213.900 1274.130 213.960 ;
        RECT 1275.190 213.900 1275.510 213.960 ;
        RECT 1273.810 172.620 1274.130 172.680 ;
        RECT 1274.270 172.620 1274.590 172.680 ;
        RECT 1273.810 172.480 1274.590 172.620 ;
        RECT 1273.810 172.420 1274.130 172.480 ;
        RECT 1274.270 172.420 1274.590 172.480 ;
        RECT 1215.850 20.300 1216.170 20.360 ;
        RECT 1274.270 20.300 1274.590 20.360 ;
        RECT 1215.850 20.160 1274.590 20.300 ;
        RECT 1215.850 20.100 1216.170 20.160 ;
        RECT 1274.270 20.100 1274.590 20.160 ;
      LAYER via ;
        RECT 1274.760 1669.440 1275.020 1669.700 ;
        RECT 1274.300 1580.360 1274.560 1580.620 ;
        RECT 1273.840 1524.600 1274.100 1524.860 ;
        RECT 1275.220 1524.600 1275.480 1524.860 ;
        RECT 1274.300 1476.320 1274.560 1476.580 ;
        RECT 1274.300 1428.380 1274.560 1428.640 ;
        RECT 1274.300 1256.000 1274.560 1256.260 ;
        RECT 1274.300 1248.860 1274.560 1249.120 ;
        RECT 1273.840 1110.820 1274.100 1111.080 ;
        RECT 1274.300 1110.480 1274.560 1110.740 ;
        RECT 1274.300 1014.260 1274.560 1014.520 ;
        RECT 1274.760 1014.260 1275.020 1014.520 ;
        RECT 1273.840 944.900 1274.100 945.160 ;
        RECT 1274.760 896.960 1275.020 897.220 ;
        RECT 1274.760 841.540 1275.020 841.800 ;
        RECT 1274.300 793.600 1274.560 793.860 ;
        RECT 1274.300 752.120 1274.560 752.380 ;
        RECT 1275.220 752.120 1275.480 752.380 ;
        RECT 1274.760 703.500 1275.020 703.760 ;
        RECT 1275.220 703.500 1275.480 703.760 ;
        RECT 1274.760 628.020 1275.020 628.280 ;
        RECT 1274.300 627.680 1274.560 627.940 ;
        RECT 1274.300 620.540 1274.560 620.800 ;
        RECT 1275.680 620.540 1275.940 620.800 ;
        RECT 1275.680 613.740 1275.940 614.000 ;
        RECT 1275.220 565.800 1275.480 566.060 ;
        RECT 1274.300 523.980 1274.560 524.240 ;
        RECT 1275.220 476.040 1275.480 476.300 ;
        RECT 1273.840 407.020 1274.100 407.280 ;
        RECT 1274.760 407.020 1275.020 407.280 ;
        RECT 1274.300 302.980 1274.560 303.240 ;
        RECT 1275.220 255.380 1275.480 255.640 ;
        RECT 1273.840 213.900 1274.100 214.160 ;
        RECT 1275.220 213.900 1275.480 214.160 ;
        RECT 1273.840 172.420 1274.100 172.680 ;
        RECT 1274.300 172.420 1274.560 172.680 ;
        RECT 1215.880 20.100 1216.140 20.360 ;
        RECT 1274.300 20.100 1274.560 20.360 ;
      LAYER met2 ;
        RECT 1274.660 1700.340 1274.940 1704.000 ;
        RECT 1274.660 1700.000 1274.960 1700.340 ;
        RECT 1274.820 1669.730 1274.960 1700.000 ;
        RECT 1274.760 1669.410 1275.020 1669.730 ;
        RECT 1274.300 1580.330 1274.560 1580.650 ;
        RECT 1274.360 1573.365 1274.500 1580.330 ;
        RECT 1274.290 1572.995 1274.570 1573.365 ;
        RECT 1273.830 1524.715 1274.110 1525.085 ;
        RECT 1273.840 1524.570 1274.100 1524.715 ;
        RECT 1275.220 1524.570 1275.480 1524.890 ;
        RECT 1275.280 1476.805 1275.420 1524.570 ;
        RECT 1274.290 1476.435 1274.570 1476.805 ;
        RECT 1275.210 1476.435 1275.490 1476.805 ;
        RECT 1274.300 1476.290 1274.560 1476.435 ;
        RECT 1274.300 1428.350 1274.560 1428.670 ;
        RECT 1274.360 1403.930 1274.500 1428.350 ;
        RECT 1274.360 1403.790 1275.420 1403.930 ;
        RECT 1275.280 1400.530 1275.420 1403.790 ;
        RECT 1274.820 1400.390 1275.420 1400.530 ;
        RECT 1274.820 1297.170 1274.960 1400.390 ;
        RECT 1274.360 1297.030 1274.960 1297.170 ;
        RECT 1274.360 1256.290 1274.500 1297.030 ;
        RECT 1274.300 1255.970 1274.560 1256.290 ;
        RECT 1274.300 1248.830 1274.560 1249.150 ;
        RECT 1274.360 1158.450 1274.500 1248.830 ;
        RECT 1273.900 1158.310 1274.500 1158.450 ;
        RECT 1273.900 1111.110 1274.040 1158.310 ;
        RECT 1273.840 1110.790 1274.100 1111.110 ;
        RECT 1274.300 1110.450 1274.560 1110.770 ;
        RECT 1274.360 1091.130 1274.500 1110.450 ;
        RECT 1274.360 1090.990 1274.960 1091.130 ;
        RECT 1274.820 1014.550 1274.960 1090.990 ;
        RECT 1274.300 1014.230 1274.560 1014.550 ;
        RECT 1274.760 1014.230 1275.020 1014.550 ;
        RECT 1274.360 946.290 1274.500 1014.230 ;
        RECT 1273.900 946.150 1274.500 946.290 ;
        RECT 1273.900 945.190 1274.040 946.150 ;
        RECT 1273.840 944.870 1274.100 945.190 ;
        RECT 1274.760 896.930 1275.020 897.250 ;
        RECT 1274.820 841.830 1274.960 896.930 ;
        RECT 1274.760 841.510 1275.020 841.830 ;
        RECT 1274.300 793.570 1274.560 793.890 ;
        RECT 1274.360 752.410 1274.500 793.570 ;
        RECT 1274.300 752.090 1274.560 752.410 ;
        RECT 1275.220 752.090 1275.480 752.410 ;
        RECT 1275.280 710.330 1275.420 752.090 ;
        RECT 1274.820 710.190 1275.420 710.330 ;
        RECT 1274.820 703.790 1274.960 710.190 ;
        RECT 1274.760 703.470 1275.020 703.790 ;
        RECT 1275.220 703.470 1275.480 703.790 ;
        RECT 1275.280 676.160 1275.420 703.470 ;
        RECT 1274.820 676.020 1275.420 676.160 ;
        RECT 1274.820 628.310 1274.960 676.020 ;
        RECT 1274.760 627.990 1275.020 628.310 ;
        RECT 1274.300 627.650 1274.560 627.970 ;
        RECT 1274.360 620.830 1274.500 627.650 ;
        RECT 1274.300 620.510 1274.560 620.830 ;
        RECT 1275.680 620.510 1275.940 620.830 ;
        RECT 1275.740 614.030 1275.880 620.510 ;
        RECT 1275.680 613.710 1275.940 614.030 ;
        RECT 1275.220 565.770 1275.480 566.090 ;
        RECT 1275.280 530.810 1275.420 565.770 ;
        RECT 1274.360 530.670 1275.420 530.810 ;
        RECT 1274.360 524.270 1274.500 530.670 ;
        RECT 1274.300 523.950 1274.560 524.270 ;
        RECT 1275.220 476.010 1275.480 476.330 ;
        RECT 1275.280 455.445 1275.420 476.010 ;
        RECT 1273.830 455.075 1274.110 455.445 ;
        RECT 1275.210 455.075 1275.490 455.445 ;
        RECT 1273.900 407.310 1274.040 455.075 ;
        RECT 1274.820 407.310 1274.960 407.465 ;
        RECT 1273.840 406.990 1274.100 407.310 ;
        RECT 1274.760 407.050 1275.020 407.310 ;
        RECT 1274.360 406.990 1275.020 407.050 ;
        RECT 1274.360 406.910 1274.960 406.990 ;
        RECT 1274.360 400.365 1274.500 406.910 ;
        RECT 1274.290 399.995 1274.570 400.365 ;
        RECT 1275.210 399.995 1275.490 400.365 ;
        RECT 1275.280 352.085 1275.420 399.995 ;
        RECT 1274.290 351.715 1274.570 352.085 ;
        RECT 1275.210 351.715 1275.490 352.085 ;
        RECT 1274.360 303.270 1274.500 351.715 ;
        RECT 1274.300 302.950 1274.560 303.270 ;
        RECT 1275.220 255.350 1275.480 255.670 ;
        RECT 1275.280 214.190 1275.420 255.350 ;
        RECT 1273.840 213.870 1274.100 214.190 ;
        RECT 1275.220 213.870 1275.480 214.190 ;
        RECT 1273.900 172.710 1274.040 213.870 ;
        RECT 1273.840 172.390 1274.100 172.710 ;
        RECT 1274.300 172.390 1274.560 172.710 ;
        RECT 1274.360 65.690 1274.500 172.390 ;
        RECT 1273.900 65.550 1274.500 65.690 ;
        RECT 1273.900 41.380 1274.040 65.550 ;
        RECT 1273.900 41.240 1274.500 41.380 ;
        RECT 1274.360 20.390 1274.500 41.240 ;
        RECT 1215.880 20.070 1216.140 20.390 ;
        RECT 1274.300 20.070 1274.560 20.390 ;
        RECT 1215.940 2.400 1216.080 20.070 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
      LAYER via2 ;
        RECT 1274.290 1573.040 1274.570 1573.320 ;
        RECT 1273.830 1524.760 1274.110 1525.040 ;
        RECT 1274.290 1476.480 1274.570 1476.760 ;
        RECT 1275.210 1476.480 1275.490 1476.760 ;
        RECT 1273.830 455.120 1274.110 455.400 ;
        RECT 1275.210 455.120 1275.490 455.400 ;
        RECT 1274.290 400.040 1274.570 400.320 ;
        RECT 1275.210 400.040 1275.490 400.320 ;
        RECT 1274.290 351.760 1274.570 352.040 ;
        RECT 1275.210 351.760 1275.490 352.040 ;
      LAYER met3 ;
        RECT 1273.550 1573.330 1273.930 1573.340 ;
        RECT 1274.265 1573.330 1274.595 1573.345 ;
        RECT 1273.550 1573.030 1274.595 1573.330 ;
        RECT 1273.550 1573.020 1273.930 1573.030 ;
        RECT 1274.265 1573.015 1274.595 1573.030 ;
        RECT 1273.805 1525.060 1274.135 1525.065 ;
        RECT 1273.550 1525.050 1274.135 1525.060 ;
        RECT 1273.550 1524.750 1274.360 1525.050 ;
        RECT 1273.550 1524.740 1274.135 1524.750 ;
        RECT 1273.805 1524.735 1274.135 1524.740 ;
        RECT 1274.265 1476.770 1274.595 1476.785 ;
        RECT 1275.185 1476.770 1275.515 1476.785 ;
        RECT 1274.265 1476.470 1275.515 1476.770 ;
        RECT 1274.265 1476.455 1274.595 1476.470 ;
        RECT 1275.185 1476.455 1275.515 1476.470 ;
        RECT 1273.805 455.410 1274.135 455.425 ;
        RECT 1275.185 455.410 1275.515 455.425 ;
        RECT 1273.805 455.110 1275.515 455.410 ;
        RECT 1273.805 455.095 1274.135 455.110 ;
        RECT 1275.185 455.095 1275.515 455.110 ;
        RECT 1274.265 400.330 1274.595 400.345 ;
        RECT 1275.185 400.330 1275.515 400.345 ;
        RECT 1274.265 400.030 1275.515 400.330 ;
        RECT 1274.265 400.015 1274.595 400.030 ;
        RECT 1275.185 400.015 1275.515 400.030 ;
        RECT 1274.265 352.050 1274.595 352.065 ;
        RECT 1275.185 352.050 1275.515 352.065 ;
        RECT 1274.265 351.750 1275.515 352.050 ;
        RECT 1274.265 351.735 1274.595 351.750 ;
        RECT 1275.185 351.735 1275.515 351.750 ;
      LAYER via3 ;
        RECT 1273.580 1573.020 1273.900 1573.340 ;
        RECT 1273.580 1524.740 1273.900 1525.060 ;
      LAYER met4 ;
        RECT 1273.575 1573.015 1273.905 1573.345 ;
        RECT 1273.590 1525.065 1273.890 1573.015 ;
        RECT 1273.575 1524.735 1273.905 1525.065 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1233.790 16.900 1234.110 16.960 ;
        RECT 1277.950 16.900 1278.270 16.960 ;
        RECT 1233.790 16.760 1278.270 16.900 ;
        RECT 1233.790 16.700 1234.110 16.760 ;
        RECT 1277.950 16.700 1278.270 16.760 ;
      LAYER via ;
        RECT 1233.820 16.700 1234.080 16.960 ;
        RECT 1277.980 16.700 1278.240 16.960 ;
      LAYER met2 ;
        RECT 1276.500 1700.340 1276.780 1704.000 ;
        RECT 1276.500 1700.000 1276.800 1700.340 ;
        RECT 1276.660 1675.930 1276.800 1700.000 ;
        RECT 1276.660 1675.790 1278.180 1675.930 ;
        RECT 1278.040 16.990 1278.180 1675.790 ;
        RECT 1233.820 16.670 1234.080 16.990 ;
        RECT 1277.980 16.670 1278.240 16.990 ;
        RECT 1233.880 2.400 1234.020 16.670 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1251.730 19.280 1252.050 19.340 ;
        RECT 1279.790 19.280 1280.110 19.340 ;
        RECT 1251.730 19.140 1280.110 19.280 ;
        RECT 1251.730 19.080 1252.050 19.140 ;
        RECT 1279.790 19.080 1280.110 19.140 ;
      LAYER via ;
        RECT 1251.760 19.080 1252.020 19.340 ;
        RECT 1279.820 19.080 1280.080 19.340 ;
      LAYER met2 ;
        RECT 1278.340 1700.340 1278.620 1704.000 ;
        RECT 1278.340 1700.000 1278.640 1700.340 ;
        RECT 1278.500 1677.290 1278.640 1700.000 ;
        RECT 1278.500 1677.150 1280.020 1677.290 ;
        RECT 1279.880 787.170 1280.020 1677.150 ;
        RECT 1279.880 787.030 1280.480 787.170 ;
        RECT 1280.340 785.130 1280.480 787.030 ;
        RECT 1279.880 784.990 1280.480 785.130 ;
        RECT 1279.880 19.370 1280.020 784.990 ;
        RECT 1251.760 19.050 1252.020 19.370 ;
        RECT 1279.820 19.050 1280.080 19.370 ;
        RECT 1251.820 2.400 1251.960 19.050 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1279.405 1642.285 1279.575 1678.495 ;
        RECT 1278.945 1445.425 1279.115 1476.535 ;
        RECT 1278.945 1324.725 1279.115 1373.175 ;
        RECT 1278.945 1187.025 1279.115 1276.275 ;
        RECT 1279.405 1041.845 1279.575 1089.955 ;
        RECT 1278.945 956.505 1279.115 993.395 ;
        RECT 1278.945 920.805 1279.115 945.115 ;
        RECT 1279.405 772.565 1279.575 787.015 ;
        RECT 1278.945 317.645 1279.115 365.415 ;
        RECT 1278.945 262.225 1279.115 309.995 ;
        RECT 1279.405 213.945 1279.575 221.255 ;
      LAYER mcon ;
        RECT 1279.405 1678.325 1279.575 1678.495 ;
        RECT 1278.945 1476.365 1279.115 1476.535 ;
        RECT 1278.945 1373.005 1279.115 1373.175 ;
        RECT 1278.945 1276.105 1279.115 1276.275 ;
        RECT 1279.405 1089.785 1279.575 1089.955 ;
        RECT 1278.945 993.225 1279.115 993.395 ;
        RECT 1278.945 944.945 1279.115 945.115 ;
        RECT 1279.405 786.845 1279.575 787.015 ;
        RECT 1278.945 365.245 1279.115 365.415 ;
        RECT 1278.945 309.825 1279.115 309.995 ;
        RECT 1279.405 221.085 1279.575 221.255 ;
      LAYER met1 ;
        RECT 1279.345 1678.480 1279.635 1678.525 ;
        RECT 1280.250 1678.480 1280.570 1678.540 ;
        RECT 1279.345 1678.340 1280.570 1678.480 ;
        RECT 1279.345 1678.295 1279.635 1678.340 ;
        RECT 1280.250 1678.280 1280.570 1678.340 ;
        RECT 1279.330 1642.440 1279.650 1642.500 ;
        RECT 1279.135 1642.300 1279.650 1642.440 ;
        RECT 1279.330 1642.240 1279.650 1642.300 ;
        RECT 1278.885 1476.520 1279.175 1476.565 ;
        RECT 1279.330 1476.520 1279.650 1476.580 ;
        RECT 1278.885 1476.380 1279.650 1476.520 ;
        RECT 1278.885 1476.335 1279.175 1476.380 ;
        RECT 1279.330 1476.320 1279.650 1476.380 ;
        RECT 1278.870 1445.580 1279.190 1445.640 ;
        RECT 1278.675 1445.440 1279.190 1445.580 ;
        RECT 1278.870 1445.380 1279.190 1445.440 ;
        RECT 1278.870 1373.160 1279.190 1373.220 ;
        RECT 1278.675 1373.020 1279.190 1373.160 ;
        RECT 1278.870 1372.960 1279.190 1373.020 ;
        RECT 1278.870 1324.880 1279.190 1324.940 ;
        RECT 1278.675 1324.740 1279.190 1324.880 ;
        RECT 1278.870 1324.680 1279.190 1324.740 ;
        RECT 1278.870 1276.260 1279.190 1276.320 ;
        RECT 1278.675 1276.120 1279.190 1276.260 ;
        RECT 1278.870 1276.060 1279.190 1276.120 ;
        RECT 1278.885 1187.180 1279.175 1187.225 ;
        RECT 1279.330 1187.180 1279.650 1187.240 ;
        RECT 1278.885 1187.040 1279.650 1187.180 ;
        RECT 1278.885 1186.995 1279.175 1187.040 ;
        RECT 1279.330 1186.980 1279.650 1187.040 ;
        RECT 1279.330 1097.760 1279.650 1097.820 ;
        RECT 1280.250 1097.760 1280.570 1097.820 ;
        RECT 1279.330 1097.620 1280.570 1097.760 ;
        RECT 1279.330 1097.560 1279.650 1097.620 ;
        RECT 1280.250 1097.560 1280.570 1097.620 ;
        RECT 1279.330 1089.940 1279.650 1090.000 ;
        RECT 1279.135 1089.800 1279.650 1089.940 ;
        RECT 1279.330 1089.740 1279.650 1089.800 ;
        RECT 1279.330 1042.000 1279.650 1042.060 ;
        RECT 1279.135 1041.860 1279.650 1042.000 ;
        RECT 1279.330 1041.800 1279.650 1041.860 ;
        RECT 1278.885 993.380 1279.175 993.425 ;
        RECT 1279.330 993.380 1279.650 993.440 ;
        RECT 1278.885 993.240 1279.650 993.380 ;
        RECT 1278.885 993.195 1279.175 993.240 ;
        RECT 1279.330 993.180 1279.650 993.240 ;
        RECT 1278.870 956.660 1279.190 956.720 ;
        RECT 1278.675 956.520 1279.190 956.660 ;
        RECT 1278.870 956.460 1279.190 956.520 ;
        RECT 1278.870 945.100 1279.190 945.160 ;
        RECT 1278.675 944.960 1279.190 945.100 ;
        RECT 1278.870 944.900 1279.190 944.960 ;
        RECT 1278.885 920.960 1279.175 921.005 ;
        RECT 1279.330 920.960 1279.650 921.020 ;
        RECT 1278.885 920.820 1279.650 920.960 ;
        RECT 1278.885 920.775 1279.175 920.820 ;
        RECT 1279.330 920.760 1279.650 920.820 ;
        RECT 1279.330 787.000 1279.650 787.060 ;
        RECT 1279.135 786.860 1279.650 787.000 ;
        RECT 1279.330 786.800 1279.650 786.860 ;
        RECT 1279.330 772.720 1279.650 772.780 ;
        RECT 1279.135 772.580 1279.650 772.720 ;
        RECT 1279.330 772.520 1279.650 772.580 ;
        RECT 1279.330 676.160 1279.650 676.220 ;
        RECT 1280.250 676.160 1280.570 676.220 ;
        RECT 1279.330 676.020 1280.570 676.160 ;
        RECT 1279.330 675.960 1279.650 676.020 ;
        RECT 1280.250 675.960 1280.570 676.020 ;
        RECT 1279.330 620.740 1279.650 620.800 ;
        RECT 1280.250 620.740 1280.570 620.800 ;
        RECT 1279.330 620.600 1280.570 620.740 ;
        RECT 1279.330 620.540 1279.650 620.600 ;
        RECT 1280.250 620.540 1280.570 620.600 ;
        RECT 1279.330 493.580 1279.650 493.640 ;
        RECT 1280.250 493.580 1280.570 493.640 ;
        RECT 1279.330 493.440 1280.570 493.580 ;
        RECT 1279.330 493.380 1279.650 493.440 ;
        RECT 1280.250 493.380 1280.570 493.440 ;
        RECT 1278.870 407.220 1279.190 407.280 ;
        RECT 1280.250 407.220 1280.570 407.280 ;
        RECT 1278.870 407.080 1280.570 407.220 ;
        RECT 1278.870 407.020 1279.190 407.080 ;
        RECT 1280.250 407.020 1280.570 407.080 ;
        RECT 1278.870 365.400 1279.190 365.460 ;
        RECT 1278.675 365.260 1279.190 365.400 ;
        RECT 1278.870 365.200 1279.190 365.260 ;
        RECT 1278.885 317.800 1279.175 317.845 ;
        RECT 1279.330 317.800 1279.650 317.860 ;
        RECT 1278.885 317.660 1279.650 317.800 ;
        RECT 1278.885 317.615 1279.175 317.660 ;
        RECT 1279.330 317.600 1279.650 317.660 ;
        RECT 1278.870 309.980 1279.190 310.040 ;
        RECT 1278.675 309.840 1279.190 309.980 ;
        RECT 1278.870 309.780 1279.190 309.840 ;
        RECT 1278.870 262.380 1279.190 262.440 ;
        RECT 1278.675 262.240 1279.190 262.380 ;
        RECT 1278.870 262.180 1279.190 262.240 ;
        RECT 1278.870 221.240 1279.190 221.300 ;
        RECT 1279.345 221.240 1279.635 221.285 ;
        RECT 1278.870 221.100 1279.635 221.240 ;
        RECT 1278.870 221.040 1279.190 221.100 ;
        RECT 1279.345 221.055 1279.635 221.100 ;
        RECT 1279.330 214.100 1279.650 214.160 ;
        RECT 1279.135 213.960 1279.650 214.100 ;
        RECT 1279.330 213.900 1279.650 213.960 ;
        RECT 1278.870 172.960 1279.190 173.020 ;
        RECT 1278.870 172.820 1279.560 172.960 ;
        RECT 1278.870 172.760 1279.190 172.820 ;
        RECT 1279.420 172.680 1279.560 172.820 ;
        RECT 1279.330 172.420 1279.650 172.680 ;
        RECT 1269.210 41.380 1269.530 41.440 ;
        RECT 1279.330 41.380 1279.650 41.440 ;
        RECT 1269.210 41.240 1279.650 41.380 ;
        RECT 1269.210 41.180 1269.530 41.240 ;
        RECT 1279.330 41.180 1279.650 41.240 ;
      LAYER via ;
        RECT 1280.280 1678.280 1280.540 1678.540 ;
        RECT 1279.360 1642.240 1279.620 1642.500 ;
        RECT 1279.360 1476.320 1279.620 1476.580 ;
        RECT 1278.900 1445.380 1279.160 1445.640 ;
        RECT 1278.900 1372.960 1279.160 1373.220 ;
        RECT 1278.900 1324.680 1279.160 1324.940 ;
        RECT 1278.900 1276.060 1279.160 1276.320 ;
        RECT 1279.360 1186.980 1279.620 1187.240 ;
        RECT 1279.360 1097.560 1279.620 1097.820 ;
        RECT 1280.280 1097.560 1280.540 1097.820 ;
        RECT 1279.360 1089.740 1279.620 1090.000 ;
        RECT 1279.360 1041.800 1279.620 1042.060 ;
        RECT 1279.360 993.180 1279.620 993.440 ;
        RECT 1278.900 956.460 1279.160 956.720 ;
        RECT 1278.900 944.900 1279.160 945.160 ;
        RECT 1279.360 920.760 1279.620 921.020 ;
        RECT 1279.360 786.800 1279.620 787.060 ;
        RECT 1279.360 772.520 1279.620 772.780 ;
        RECT 1279.360 675.960 1279.620 676.220 ;
        RECT 1280.280 675.960 1280.540 676.220 ;
        RECT 1279.360 620.540 1279.620 620.800 ;
        RECT 1280.280 620.540 1280.540 620.800 ;
        RECT 1279.360 493.380 1279.620 493.640 ;
        RECT 1280.280 493.380 1280.540 493.640 ;
        RECT 1278.900 407.020 1279.160 407.280 ;
        RECT 1280.280 407.020 1280.540 407.280 ;
        RECT 1278.900 365.200 1279.160 365.460 ;
        RECT 1279.360 317.600 1279.620 317.860 ;
        RECT 1278.900 309.780 1279.160 310.040 ;
        RECT 1278.900 262.180 1279.160 262.440 ;
        RECT 1278.900 221.040 1279.160 221.300 ;
        RECT 1279.360 213.900 1279.620 214.160 ;
        RECT 1278.900 172.760 1279.160 173.020 ;
        RECT 1279.360 172.420 1279.620 172.680 ;
        RECT 1269.240 41.180 1269.500 41.440 ;
        RECT 1279.360 41.180 1279.620 41.440 ;
      LAYER met2 ;
        RECT 1280.180 1700.340 1280.460 1704.000 ;
        RECT 1280.180 1700.000 1280.480 1700.340 ;
        RECT 1280.340 1678.570 1280.480 1700.000 ;
        RECT 1280.280 1678.250 1280.540 1678.570 ;
        RECT 1279.360 1642.210 1279.620 1642.530 ;
        RECT 1279.420 1486.890 1279.560 1642.210 ;
        RECT 1278.960 1486.750 1279.560 1486.890 ;
        RECT 1278.960 1483.490 1279.100 1486.750 ;
        RECT 1278.960 1483.350 1279.560 1483.490 ;
        RECT 1279.420 1476.610 1279.560 1483.350 ;
        RECT 1279.360 1476.290 1279.620 1476.610 ;
        RECT 1278.900 1445.525 1279.160 1445.670 ;
        RECT 1278.890 1445.155 1279.170 1445.525 ;
        RECT 1278.890 1379.875 1279.170 1380.245 ;
        RECT 1278.960 1373.250 1279.100 1379.875 ;
        RECT 1278.900 1372.930 1279.160 1373.250 ;
        RECT 1278.900 1324.650 1279.160 1324.970 ;
        RECT 1278.960 1276.350 1279.100 1324.650 ;
        RECT 1278.900 1276.030 1279.160 1276.350 ;
        RECT 1279.360 1186.950 1279.620 1187.270 ;
        RECT 1279.420 1186.330 1279.560 1186.950 ;
        RECT 1278.960 1186.190 1279.560 1186.330 ;
        RECT 1278.960 1138.845 1279.100 1186.190 ;
        RECT 1278.890 1138.475 1279.170 1138.845 ;
        RECT 1280.270 1138.475 1280.550 1138.845 ;
        RECT 1280.340 1097.850 1280.480 1138.475 ;
        RECT 1279.360 1097.530 1279.620 1097.850 ;
        RECT 1280.280 1097.530 1280.540 1097.850 ;
        RECT 1279.420 1090.030 1279.560 1097.530 ;
        RECT 1279.360 1089.710 1279.620 1090.030 ;
        RECT 1279.360 1041.770 1279.620 1042.090 ;
        RECT 1279.420 993.470 1279.560 1041.770 ;
        RECT 1279.360 993.150 1279.620 993.470 ;
        RECT 1278.900 956.430 1279.160 956.750 ;
        RECT 1278.960 945.190 1279.100 956.430 ;
        RECT 1278.900 944.870 1279.160 945.190 ;
        RECT 1279.360 920.730 1279.620 921.050 ;
        RECT 1279.420 787.090 1279.560 920.730 ;
        RECT 1279.360 786.770 1279.620 787.090 ;
        RECT 1279.360 772.490 1279.620 772.810 ;
        RECT 1279.420 676.250 1279.560 772.490 ;
        RECT 1279.360 675.930 1279.620 676.250 ;
        RECT 1280.280 675.930 1280.540 676.250 ;
        RECT 1280.340 628.165 1280.480 675.930 ;
        RECT 1279.350 627.795 1279.630 628.165 ;
        RECT 1280.270 627.795 1280.550 628.165 ;
        RECT 1279.420 620.830 1279.560 627.795 ;
        RECT 1279.360 620.510 1279.620 620.830 ;
        RECT 1280.280 620.510 1280.540 620.830 ;
        RECT 1280.340 531.605 1280.480 620.510 ;
        RECT 1279.350 531.235 1279.630 531.605 ;
        RECT 1280.270 531.235 1280.550 531.605 ;
        RECT 1279.420 493.670 1279.560 531.235 ;
        RECT 1279.360 493.350 1279.620 493.670 ;
        RECT 1280.280 493.350 1280.540 493.670 ;
        RECT 1280.340 407.310 1280.480 493.350 ;
        RECT 1278.900 406.990 1279.160 407.310 ;
        RECT 1280.280 406.990 1280.540 407.310 ;
        RECT 1278.960 365.490 1279.100 406.990 ;
        RECT 1278.900 365.170 1279.160 365.490 ;
        RECT 1279.360 317.570 1279.620 317.890 ;
        RECT 1279.420 310.490 1279.560 317.570 ;
        RECT 1278.960 310.350 1279.560 310.490 ;
        RECT 1278.960 310.070 1279.100 310.350 ;
        RECT 1278.900 309.750 1279.160 310.070 ;
        RECT 1278.900 262.150 1279.160 262.470 ;
        RECT 1278.960 221.330 1279.100 262.150 ;
        RECT 1278.900 221.010 1279.160 221.330 ;
        RECT 1279.360 214.100 1279.620 214.190 ;
        RECT 1278.960 213.960 1279.620 214.100 ;
        RECT 1278.960 173.050 1279.100 213.960 ;
        RECT 1279.360 213.870 1279.620 213.960 ;
        RECT 1278.900 172.730 1279.160 173.050 ;
        RECT 1279.360 172.390 1279.620 172.710 ;
        RECT 1279.420 41.470 1279.560 172.390 ;
        RECT 1269.240 41.150 1269.500 41.470 ;
        RECT 1279.360 41.150 1279.620 41.470 ;
        RECT 1269.300 2.400 1269.440 41.150 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
      LAYER via2 ;
        RECT 1278.890 1445.200 1279.170 1445.480 ;
        RECT 1278.890 1379.920 1279.170 1380.200 ;
        RECT 1278.890 1138.520 1279.170 1138.800 ;
        RECT 1280.270 1138.520 1280.550 1138.800 ;
        RECT 1279.350 627.840 1279.630 628.120 ;
        RECT 1280.270 627.840 1280.550 628.120 ;
        RECT 1279.350 531.280 1279.630 531.560 ;
        RECT 1280.270 531.280 1280.550 531.560 ;
      LAYER met3 ;
        RECT 1278.150 1445.490 1278.530 1445.500 ;
        RECT 1278.865 1445.490 1279.195 1445.505 ;
        RECT 1278.150 1445.190 1279.195 1445.490 ;
        RECT 1278.150 1445.180 1278.530 1445.190 ;
        RECT 1278.865 1445.175 1279.195 1445.190 ;
        RECT 1278.150 1380.210 1278.530 1380.220 ;
        RECT 1278.865 1380.210 1279.195 1380.225 ;
        RECT 1278.150 1379.910 1279.195 1380.210 ;
        RECT 1278.150 1379.900 1278.530 1379.910 ;
        RECT 1278.865 1379.895 1279.195 1379.910 ;
        RECT 1278.865 1138.810 1279.195 1138.825 ;
        RECT 1280.245 1138.810 1280.575 1138.825 ;
        RECT 1278.865 1138.510 1280.575 1138.810 ;
        RECT 1278.865 1138.495 1279.195 1138.510 ;
        RECT 1280.245 1138.495 1280.575 1138.510 ;
        RECT 1279.325 628.130 1279.655 628.145 ;
        RECT 1280.245 628.130 1280.575 628.145 ;
        RECT 1279.325 627.830 1280.575 628.130 ;
        RECT 1279.325 627.815 1279.655 627.830 ;
        RECT 1280.245 627.815 1280.575 627.830 ;
        RECT 1279.325 531.570 1279.655 531.585 ;
        RECT 1280.245 531.570 1280.575 531.585 ;
        RECT 1279.325 531.270 1280.575 531.570 ;
        RECT 1279.325 531.255 1279.655 531.270 ;
        RECT 1280.245 531.255 1280.575 531.270 ;
      LAYER via3 ;
        RECT 1278.180 1445.180 1278.500 1445.500 ;
        RECT 1278.180 1379.900 1278.500 1380.220 ;
      LAYER met4 ;
        RECT 1278.175 1445.175 1278.505 1445.505 ;
        RECT 1278.190 1380.225 1278.490 1445.175 ;
        RECT 1278.175 1379.895 1278.505 1380.225 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1282.625 476.085 1282.795 524.195 ;
        RECT 1282.165 317.645 1282.335 365.755 ;
        RECT 1283.085 89.845 1283.255 220.575 ;
        RECT 1282.625 41.565 1282.795 48.535 ;
      LAYER mcon ;
        RECT 1282.625 524.025 1282.795 524.195 ;
        RECT 1282.165 365.585 1282.335 365.755 ;
        RECT 1283.085 220.405 1283.255 220.575 ;
        RECT 1282.625 48.365 1282.795 48.535 ;
      LAYER met1 ;
        RECT 1282.090 1640.740 1282.410 1640.800 ;
        RECT 1283.470 1640.740 1283.790 1640.800 ;
        RECT 1282.090 1640.600 1283.790 1640.740 ;
        RECT 1282.090 1640.540 1282.410 1640.600 ;
        RECT 1283.470 1640.540 1283.790 1640.600 ;
        RECT 1283.010 1580.560 1283.330 1580.620 ;
        RECT 1283.470 1580.560 1283.790 1580.620 ;
        RECT 1283.010 1580.420 1283.790 1580.560 ;
        RECT 1283.010 1580.360 1283.330 1580.420 ;
        RECT 1283.470 1580.360 1283.790 1580.420 ;
        RECT 1282.090 1476.520 1282.410 1476.580 ;
        RECT 1283.010 1476.520 1283.330 1476.580 ;
        RECT 1282.090 1476.380 1283.330 1476.520 ;
        RECT 1282.090 1476.320 1282.410 1476.380 ;
        RECT 1283.010 1476.320 1283.330 1476.380 ;
        RECT 1282.550 1193.640 1282.870 1193.700 ;
        RECT 1283.010 1193.640 1283.330 1193.700 ;
        RECT 1282.550 1193.500 1283.330 1193.640 ;
        RECT 1282.550 1193.440 1282.870 1193.500 ;
        RECT 1283.010 1193.440 1283.330 1193.500 ;
        RECT 1283.010 1104.560 1283.330 1104.620 ;
        RECT 1282.180 1104.420 1283.330 1104.560 ;
        RECT 1282.180 1103.940 1282.320 1104.420 ;
        RECT 1283.010 1104.360 1283.330 1104.420 ;
        RECT 1282.090 1103.680 1282.410 1103.940 ;
        RECT 1282.550 524.180 1282.870 524.240 ;
        RECT 1282.355 524.040 1282.870 524.180 ;
        RECT 1282.550 523.980 1282.870 524.040 ;
        RECT 1282.565 476.240 1282.855 476.285 ;
        RECT 1283.470 476.240 1283.790 476.300 ;
        RECT 1282.565 476.100 1283.790 476.240 ;
        RECT 1282.565 476.055 1282.855 476.100 ;
        RECT 1283.470 476.040 1283.790 476.100 ;
        RECT 1282.090 414.020 1282.410 414.080 ;
        RECT 1283.010 414.020 1283.330 414.080 ;
        RECT 1282.090 413.880 1283.330 414.020 ;
        RECT 1282.090 413.820 1282.410 413.880 ;
        RECT 1283.010 413.820 1283.330 413.880 ;
        RECT 1282.090 365.740 1282.410 365.800 ;
        RECT 1281.895 365.600 1282.410 365.740 ;
        RECT 1282.090 365.540 1282.410 365.600 ;
        RECT 1282.105 317.800 1282.395 317.845 ;
        RECT 1283.010 317.800 1283.330 317.860 ;
        RECT 1282.105 317.660 1283.330 317.800 ;
        RECT 1282.105 317.615 1282.395 317.660 ;
        RECT 1283.010 317.600 1283.330 317.660 ;
        RECT 1283.010 220.560 1283.330 220.620 ;
        RECT 1282.815 220.420 1283.330 220.560 ;
        RECT 1283.010 220.360 1283.330 220.420 ;
        RECT 1283.010 90.000 1283.330 90.060 ;
        RECT 1282.815 89.860 1283.330 90.000 ;
        RECT 1283.010 89.800 1283.330 89.860 ;
        RECT 1282.550 48.520 1282.870 48.580 ;
        RECT 1282.355 48.380 1282.870 48.520 ;
        RECT 1282.550 48.320 1282.870 48.380 ;
        RECT 1282.550 41.720 1282.870 41.780 ;
        RECT 1282.355 41.580 1282.870 41.720 ;
        RECT 1282.550 41.520 1282.870 41.580 ;
        RECT 1282.550 9.420 1282.870 9.480 ;
        RECT 1287.150 9.420 1287.470 9.480 ;
        RECT 1282.550 9.280 1287.470 9.420 ;
        RECT 1282.550 9.220 1282.870 9.280 ;
        RECT 1287.150 9.220 1287.470 9.280 ;
      LAYER via ;
        RECT 1282.120 1640.540 1282.380 1640.800 ;
        RECT 1283.500 1640.540 1283.760 1640.800 ;
        RECT 1283.040 1580.360 1283.300 1580.620 ;
        RECT 1283.500 1580.360 1283.760 1580.620 ;
        RECT 1282.120 1476.320 1282.380 1476.580 ;
        RECT 1283.040 1476.320 1283.300 1476.580 ;
        RECT 1282.580 1193.440 1282.840 1193.700 ;
        RECT 1283.040 1193.440 1283.300 1193.700 ;
        RECT 1283.040 1104.360 1283.300 1104.620 ;
        RECT 1282.120 1103.680 1282.380 1103.940 ;
        RECT 1282.580 523.980 1282.840 524.240 ;
        RECT 1283.500 476.040 1283.760 476.300 ;
        RECT 1282.120 413.820 1282.380 414.080 ;
        RECT 1283.040 413.820 1283.300 414.080 ;
        RECT 1282.120 365.540 1282.380 365.800 ;
        RECT 1283.040 317.600 1283.300 317.860 ;
        RECT 1283.040 220.360 1283.300 220.620 ;
        RECT 1283.040 89.800 1283.300 90.060 ;
        RECT 1282.580 48.320 1282.840 48.580 ;
        RECT 1282.580 41.520 1282.840 41.780 ;
        RECT 1282.580 9.220 1282.840 9.480 ;
        RECT 1287.180 9.220 1287.440 9.480 ;
      LAYER met2 ;
        RECT 1282.020 1700.340 1282.300 1704.000 ;
        RECT 1282.020 1700.000 1282.320 1700.340 ;
        RECT 1282.180 1640.830 1282.320 1700.000 ;
        RECT 1282.120 1640.510 1282.380 1640.830 ;
        RECT 1283.500 1640.510 1283.760 1640.830 ;
        RECT 1283.560 1580.650 1283.700 1640.510 ;
        RECT 1283.040 1580.330 1283.300 1580.650 ;
        RECT 1283.500 1580.330 1283.760 1580.650 ;
        RECT 1283.100 1573.365 1283.240 1580.330 ;
        RECT 1282.110 1572.995 1282.390 1573.365 ;
        RECT 1283.030 1572.995 1283.310 1573.365 ;
        RECT 1282.180 1525.085 1282.320 1572.995 ;
        RECT 1282.110 1524.715 1282.390 1525.085 ;
        RECT 1283.030 1524.715 1283.310 1525.085 ;
        RECT 1283.100 1476.610 1283.240 1524.715 ;
        RECT 1282.120 1476.290 1282.380 1476.610 ;
        RECT 1283.040 1476.290 1283.300 1476.610 ;
        RECT 1282.180 1428.525 1282.320 1476.290 ;
        RECT 1282.110 1428.155 1282.390 1428.525 ;
        RECT 1283.030 1428.155 1283.310 1428.525 ;
        RECT 1283.100 1193.810 1283.240 1428.155 ;
        RECT 1282.640 1193.730 1283.240 1193.810 ;
        RECT 1282.580 1193.670 1283.300 1193.730 ;
        RECT 1282.580 1193.410 1282.840 1193.670 ;
        RECT 1283.040 1193.410 1283.300 1193.670 ;
        RECT 1283.100 1104.650 1283.240 1193.410 ;
        RECT 1283.040 1104.330 1283.300 1104.650 ;
        RECT 1282.120 1103.650 1282.380 1103.970 ;
        RECT 1282.180 966.125 1282.320 1103.650 ;
        RECT 1282.110 965.755 1282.390 966.125 ;
        RECT 1283.030 965.755 1283.310 966.125 ;
        RECT 1283.100 531.490 1283.240 965.755 ;
        RECT 1282.640 531.350 1283.240 531.490 ;
        RECT 1282.640 524.270 1282.780 531.350 ;
        RECT 1282.580 523.950 1282.840 524.270 ;
        RECT 1283.500 476.010 1283.760 476.330 ;
        RECT 1283.560 445.130 1283.700 476.010 ;
        RECT 1283.100 444.990 1283.700 445.130 ;
        RECT 1283.100 414.110 1283.240 444.990 ;
        RECT 1282.120 413.790 1282.380 414.110 ;
        RECT 1283.040 413.790 1283.300 414.110 ;
        RECT 1282.180 365.830 1282.320 413.790 ;
        RECT 1282.120 365.510 1282.380 365.830 ;
        RECT 1283.040 317.570 1283.300 317.890 ;
        RECT 1283.100 220.650 1283.240 317.570 ;
        RECT 1283.040 220.330 1283.300 220.650 ;
        RECT 1283.040 89.770 1283.300 90.090 ;
        RECT 1283.100 89.490 1283.240 89.770 ;
        RECT 1282.640 89.350 1283.240 89.490 ;
        RECT 1282.640 48.610 1282.780 89.350 ;
        RECT 1282.580 48.290 1282.840 48.610 ;
        RECT 1282.580 41.490 1282.840 41.810 ;
        RECT 1282.640 9.510 1282.780 41.490 ;
        RECT 1282.580 9.190 1282.840 9.510 ;
        RECT 1287.180 9.190 1287.440 9.510 ;
        RECT 1287.240 2.400 1287.380 9.190 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
      LAYER via2 ;
        RECT 1282.110 1573.040 1282.390 1573.320 ;
        RECT 1283.030 1573.040 1283.310 1573.320 ;
        RECT 1282.110 1524.760 1282.390 1525.040 ;
        RECT 1283.030 1524.760 1283.310 1525.040 ;
        RECT 1282.110 1428.200 1282.390 1428.480 ;
        RECT 1283.030 1428.200 1283.310 1428.480 ;
        RECT 1282.110 965.800 1282.390 966.080 ;
        RECT 1283.030 965.800 1283.310 966.080 ;
      LAYER met3 ;
        RECT 1282.085 1573.330 1282.415 1573.345 ;
        RECT 1283.005 1573.330 1283.335 1573.345 ;
        RECT 1282.085 1573.030 1283.335 1573.330 ;
        RECT 1282.085 1573.015 1282.415 1573.030 ;
        RECT 1283.005 1573.015 1283.335 1573.030 ;
        RECT 1282.085 1525.050 1282.415 1525.065 ;
        RECT 1283.005 1525.050 1283.335 1525.065 ;
        RECT 1282.085 1524.750 1283.335 1525.050 ;
        RECT 1282.085 1524.735 1282.415 1524.750 ;
        RECT 1283.005 1524.735 1283.335 1524.750 ;
        RECT 1282.085 1428.490 1282.415 1428.505 ;
        RECT 1283.005 1428.490 1283.335 1428.505 ;
        RECT 1282.085 1428.190 1283.335 1428.490 ;
        RECT 1282.085 1428.175 1282.415 1428.190 ;
        RECT 1283.005 1428.175 1283.335 1428.190 ;
        RECT 1282.085 966.090 1282.415 966.105 ;
        RECT 1283.005 966.090 1283.335 966.105 ;
        RECT 1282.085 965.790 1283.335 966.090 ;
        RECT 1282.085 965.775 1282.415 965.790 ;
        RECT 1283.005 965.775 1283.335 965.790 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1283.930 1684.600 1284.250 1684.660 ;
        RECT 1288.530 1684.600 1288.850 1684.660 ;
        RECT 1283.930 1684.460 1288.850 1684.600 ;
        RECT 1283.930 1684.400 1284.250 1684.460 ;
        RECT 1288.530 1684.400 1288.850 1684.460 ;
        RECT 1288.530 19.960 1288.850 20.020 ;
        RECT 1305.090 19.960 1305.410 20.020 ;
        RECT 1288.530 19.820 1305.410 19.960 ;
        RECT 1288.530 19.760 1288.850 19.820 ;
        RECT 1305.090 19.760 1305.410 19.820 ;
      LAYER via ;
        RECT 1283.960 1684.400 1284.220 1684.660 ;
        RECT 1288.560 1684.400 1288.820 1684.660 ;
        RECT 1288.560 19.760 1288.820 20.020 ;
        RECT 1305.120 19.760 1305.380 20.020 ;
      LAYER met2 ;
        RECT 1283.860 1700.340 1284.140 1704.000 ;
        RECT 1283.860 1700.000 1284.160 1700.340 ;
        RECT 1284.020 1684.690 1284.160 1700.000 ;
        RECT 1283.960 1684.370 1284.220 1684.690 ;
        RECT 1288.560 1684.370 1288.820 1684.690 ;
        RECT 1288.620 20.050 1288.760 1684.370 ;
        RECT 1288.560 19.730 1288.820 20.050 ;
        RECT 1305.120 19.730 1305.380 20.050 ;
        RECT 1305.180 2.400 1305.320 19.730 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1312.525 1681.385 1312.695 1688.015 ;
      LAYER mcon ;
        RECT 1312.525 1687.845 1312.695 1688.015 ;
      LAYER met1 ;
        RECT 1285.770 1688.000 1286.090 1688.060 ;
        RECT 1312.465 1688.000 1312.755 1688.045 ;
        RECT 1285.770 1687.860 1312.755 1688.000 ;
        RECT 1285.770 1687.800 1286.090 1687.860 ;
        RECT 1312.465 1687.815 1312.755 1687.860 ;
        RECT 1312.450 1681.540 1312.770 1681.600 ;
        RECT 1312.255 1681.400 1312.770 1681.540 ;
        RECT 1312.450 1681.340 1312.770 1681.400 ;
        RECT 1312.450 1667.260 1312.770 1667.320 ;
        RECT 1314.290 1667.260 1314.610 1667.320 ;
        RECT 1312.450 1667.120 1314.610 1667.260 ;
        RECT 1312.450 1667.060 1312.770 1667.120 ;
        RECT 1314.290 1667.060 1314.610 1667.120 ;
        RECT 1314.290 20.640 1314.610 20.700 ;
        RECT 1323.030 20.640 1323.350 20.700 ;
        RECT 1314.290 20.500 1323.350 20.640 ;
        RECT 1314.290 20.440 1314.610 20.500 ;
        RECT 1323.030 20.440 1323.350 20.500 ;
      LAYER via ;
        RECT 1285.800 1687.800 1286.060 1688.060 ;
        RECT 1312.480 1681.340 1312.740 1681.600 ;
        RECT 1312.480 1667.060 1312.740 1667.320 ;
        RECT 1314.320 1667.060 1314.580 1667.320 ;
        RECT 1314.320 20.440 1314.580 20.700 ;
        RECT 1323.060 20.440 1323.320 20.700 ;
      LAYER met2 ;
        RECT 1285.700 1700.340 1285.980 1704.000 ;
        RECT 1285.700 1700.000 1286.000 1700.340 ;
        RECT 1285.860 1688.090 1286.000 1700.000 ;
        RECT 1285.800 1687.770 1286.060 1688.090 ;
        RECT 1312.480 1681.310 1312.740 1681.630 ;
        RECT 1312.540 1667.350 1312.680 1681.310 ;
        RECT 1312.480 1667.030 1312.740 1667.350 ;
        RECT 1314.320 1667.030 1314.580 1667.350 ;
        RECT 1314.380 20.730 1314.520 1667.030 ;
        RECT 1314.320 20.410 1314.580 20.730 ;
        RECT 1323.060 20.410 1323.320 20.730 ;
        RECT 1323.120 2.400 1323.260 20.410 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1314.365 1683.425 1314.535 1687.675 ;
      LAYER mcon ;
        RECT 1314.365 1687.505 1314.535 1687.675 ;
      LAYER met1 ;
        RECT 1287.610 1687.660 1287.930 1687.720 ;
        RECT 1314.305 1687.660 1314.595 1687.705 ;
        RECT 1287.610 1687.520 1314.595 1687.660 ;
        RECT 1287.610 1687.460 1287.930 1687.520 ;
        RECT 1314.305 1687.475 1314.595 1687.520 ;
        RECT 1314.290 1683.580 1314.610 1683.640 ;
        RECT 1314.095 1683.440 1314.610 1683.580 ;
        RECT 1314.290 1683.380 1314.610 1683.440 ;
        RECT 1314.750 34.580 1315.070 34.640 ;
        RECT 1340.510 34.580 1340.830 34.640 ;
        RECT 1314.750 34.440 1340.830 34.580 ;
        RECT 1314.750 34.380 1315.070 34.440 ;
        RECT 1340.510 34.380 1340.830 34.440 ;
      LAYER via ;
        RECT 1287.640 1687.460 1287.900 1687.720 ;
        RECT 1314.320 1683.380 1314.580 1683.640 ;
        RECT 1314.780 34.380 1315.040 34.640 ;
        RECT 1340.540 34.380 1340.800 34.640 ;
      LAYER met2 ;
        RECT 1287.540 1700.340 1287.820 1704.000 ;
        RECT 1287.540 1700.000 1287.840 1700.340 ;
        RECT 1287.700 1687.750 1287.840 1700.000 ;
        RECT 1287.640 1687.430 1287.900 1687.750 ;
        RECT 1314.320 1683.350 1314.580 1683.670 ;
        RECT 1314.380 1667.770 1314.520 1683.350 ;
        RECT 1314.380 1667.630 1314.980 1667.770 ;
        RECT 1314.840 34.670 1314.980 1667.630 ;
        RECT 1314.780 34.350 1315.040 34.670 ;
        RECT 1340.540 34.350 1340.800 34.670 ;
        RECT 1340.600 2.400 1340.740 34.350 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 703.410 1583.960 703.730 1584.020 ;
        RECT 1222.750 1583.960 1223.070 1584.020 ;
        RECT 703.410 1583.820 1223.070 1583.960 ;
        RECT 703.410 1583.760 703.730 1583.820 ;
        RECT 1222.750 1583.760 1223.070 1583.820 ;
      LAYER via ;
        RECT 703.440 1583.760 703.700 1584.020 ;
        RECT 1222.780 1583.760 1223.040 1584.020 ;
      LAYER met2 ;
        RECT 1221.300 1700.410 1221.580 1704.000 ;
        RECT 1221.300 1700.270 1222.060 1700.410 ;
        RECT 1221.300 1700.000 1221.580 1700.270 ;
        RECT 1221.920 1663.690 1222.060 1700.270 ;
        RECT 1221.920 1663.550 1222.980 1663.690 ;
        RECT 1222.840 1584.050 1222.980 1663.550 ;
        RECT 703.440 1583.730 703.700 1584.050 ;
        RECT 1222.780 1583.730 1223.040 1584.050 ;
        RECT 703.500 24.210 703.640 1583.730 ;
        RECT 698.440 24.070 703.640 24.210 ;
        RECT 698.440 2.400 698.580 24.070 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1287.150 1683.920 1287.470 1683.980 ;
        RECT 1289.450 1683.920 1289.770 1683.980 ;
        RECT 1287.150 1683.780 1289.770 1683.920 ;
        RECT 1287.150 1683.720 1287.470 1683.780 ;
        RECT 1289.450 1683.720 1289.770 1683.780 ;
        RECT 1287.150 1590.420 1287.470 1590.480 ;
        RECT 1352.470 1590.420 1352.790 1590.480 ;
        RECT 1287.150 1590.280 1352.790 1590.420 ;
        RECT 1287.150 1590.220 1287.470 1590.280 ;
        RECT 1352.470 1590.220 1352.790 1590.280 ;
        RECT 1352.470 7.040 1352.790 7.100 ;
        RECT 1358.450 7.040 1358.770 7.100 ;
        RECT 1352.470 6.900 1358.770 7.040 ;
        RECT 1352.470 6.840 1352.790 6.900 ;
        RECT 1358.450 6.840 1358.770 6.900 ;
      LAYER via ;
        RECT 1287.180 1683.720 1287.440 1683.980 ;
        RECT 1289.480 1683.720 1289.740 1683.980 ;
        RECT 1287.180 1590.220 1287.440 1590.480 ;
        RECT 1352.500 1590.220 1352.760 1590.480 ;
        RECT 1352.500 6.840 1352.760 7.100 ;
        RECT 1358.480 6.840 1358.740 7.100 ;
      LAYER met2 ;
        RECT 1289.380 1700.340 1289.660 1704.000 ;
        RECT 1289.380 1700.000 1289.680 1700.340 ;
        RECT 1289.540 1684.010 1289.680 1700.000 ;
        RECT 1287.180 1683.690 1287.440 1684.010 ;
        RECT 1289.480 1683.690 1289.740 1684.010 ;
        RECT 1287.240 1590.510 1287.380 1683.690 ;
        RECT 1287.180 1590.190 1287.440 1590.510 ;
        RECT 1352.500 1590.190 1352.760 1590.510 ;
        RECT 1352.560 7.130 1352.700 1590.190 ;
        RECT 1352.500 6.810 1352.760 7.130 ;
        RECT 1358.480 6.810 1358.740 7.130 ;
        RECT 1358.540 2.400 1358.680 6.810 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1362.665 1677.305 1362.835 1688.355 ;
      LAYER mcon ;
        RECT 1362.665 1688.185 1362.835 1688.355 ;
      LAYER met1 ;
        RECT 1291.290 1688.340 1291.610 1688.400 ;
        RECT 1362.605 1688.340 1362.895 1688.385 ;
        RECT 1291.290 1688.200 1362.895 1688.340 ;
        RECT 1291.290 1688.140 1291.610 1688.200 ;
        RECT 1362.605 1688.155 1362.895 1688.200 ;
        RECT 1362.590 1677.460 1362.910 1677.520 ;
        RECT 1362.395 1677.320 1362.910 1677.460 ;
        RECT 1362.590 1677.260 1362.910 1677.320 ;
        RECT 1362.590 41.380 1362.910 41.440 ;
        RECT 1376.390 41.380 1376.710 41.440 ;
        RECT 1362.590 41.240 1376.710 41.380 ;
        RECT 1362.590 41.180 1362.910 41.240 ;
        RECT 1376.390 41.180 1376.710 41.240 ;
      LAYER via ;
        RECT 1291.320 1688.140 1291.580 1688.400 ;
        RECT 1362.620 1677.260 1362.880 1677.520 ;
        RECT 1362.620 41.180 1362.880 41.440 ;
        RECT 1376.420 41.180 1376.680 41.440 ;
      LAYER met2 ;
        RECT 1291.220 1700.340 1291.500 1704.000 ;
        RECT 1291.220 1700.000 1291.520 1700.340 ;
        RECT 1291.380 1688.430 1291.520 1700.000 ;
        RECT 1291.320 1688.110 1291.580 1688.430 ;
        RECT 1362.620 1677.230 1362.880 1677.550 ;
        RECT 1362.680 41.470 1362.820 1677.230 ;
        RECT 1362.620 41.150 1362.880 41.470 ;
        RECT 1376.420 41.150 1376.680 41.470 ;
        RECT 1376.480 2.400 1376.620 41.150 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1308.845 1642.285 1309.015 1686.655 ;
      LAYER mcon ;
        RECT 1308.845 1686.485 1309.015 1686.655 ;
      LAYER met1 ;
        RECT 1293.130 1686.640 1293.450 1686.700 ;
        RECT 1308.785 1686.640 1309.075 1686.685 ;
        RECT 1293.130 1686.500 1309.075 1686.640 ;
        RECT 1293.130 1686.440 1293.450 1686.500 ;
        RECT 1308.785 1686.455 1309.075 1686.500 ;
        RECT 1308.770 1642.440 1309.090 1642.500 ;
        RECT 1308.575 1642.300 1309.090 1642.440 ;
        RECT 1308.770 1642.240 1309.090 1642.300 ;
        RECT 1308.770 1569.680 1309.090 1569.740 ;
        RECT 1393.870 1569.680 1394.190 1569.740 ;
        RECT 1308.770 1569.540 1394.190 1569.680 ;
        RECT 1308.770 1569.480 1309.090 1569.540 ;
        RECT 1393.870 1569.480 1394.190 1569.540 ;
      LAYER via ;
        RECT 1293.160 1686.440 1293.420 1686.700 ;
        RECT 1308.800 1642.240 1309.060 1642.500 ;
        RECT 1308.800 1569.480 1309.060 1569.740 ;
        RECT 1393.900 1569.480 1394.160 1569.740 ;
      LAYER met2 ;
        RECT 1293.060 1700.340 1293.340 1704.000 ;
        RECT 1293.060 1700.000 1293.360 1700.340 ;
        RECT 1293.220 1686.730 1293.360 1700.000 ;
        RECT 1293.160 1686.410 1293.420 1686.730 ;
        RECT 1308.800 1642.210 1309.060 1642.530 ;
        RECT 1308.860 1569.770 1309.000 1642.210 ;
        RECT 1308.800 1569.450 1309.060 1569.770 ;
        RECT 1393.900 1569.450 1394.160 1569.770 ;
        RECT 1393.960 3.130 1394.100 1569.450 ;
        RECT 1393.960 2.990 1394.560 3.130 ;
        RECT 1394.420 2.400 1394.560 2.990 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1294.970 1638.700 1295.290 1638.760 ;
        RECT 1407.670 1638.700 1407.990 1638.760 ;
        RECT 1294.970 1638.560 1407.990 1638.700 ;
        RECT 1294.970 1638.500 1295.290 1638.560 ;
        RECT 1407.670 1638.500 1407.990 1638.560 ;
        RECT 1407.670 2.960 1407.990 3.020 ;
        RECT 1412.270 2.960 1412.590 3.020 ;
        RECT 1407.670 2.820 1412.590 2.960 ;
        RECT 1407.670 2.760 1407.990 2.820 ;
        RECT 1412.270 2.760 1412.590 2.820 ;
      LAYER via ;
        RECT 1295.000 1638.500 1295.260 1638.760 ;
        RECT 1407.700 1638.500 1407.960 1638.760 ;
        RECT 1407.700 2.760 1407.960 3.020 ;
        RECT 1412.300 2.760 1412.560 3.020 ;
      LAYER met2 ;
        RECT 1294.900 1700.340 1295.180 1704.000 ;
        RECT 1294.900 1700.000 1295.200 1700.340 ;
        RECT 1295.060 1638.790 1295.200 1700.000 ;
        RECT 1295.000 1638.470 1295.260 1638.790 ;
        RECT 1407.700 1638.470 1407.960 1638.790 ;
        RECT 1407.760 3.050 1407.900 1638.470 ;
        RECT 1407.700 2.730 1407.960 3.050 ;
        RECT 1412.300 2.730 1412.560 3.050 ;
        RECT 1412.360 2.400 1412.500 2.730 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1291.290 1656.040 1291.610 1656.100 ;
        RECT 1296.810 1656.040 1297.130 1656.100 ;
        RECT 1291.290 1655.900 1297.130 1656.040 ;
        RECT 1291.290 1655.840 1291.610 1655.900 ;
        RECT 1296.810 1655.840 1297.130 1655.900 ;
        RECT 1291.290 1577.500 1291.610 1577.560 ;
        RECT 1428.370 1577.500 1428.690 1577.560 ;
        RECT 1291.290 1577.360 1428.690 1577.500 ;
        RECT 1291.290 1577.300 1291.610 1577.360 ;
        RECT 1428.370 1577.300 1428.690 1577.360 ;
        RECT 1428.370 2.960 1428.690 3.020 ;
        RECT 1429.750 2.960 1430.070 3.020 ;
        RECT 1428.370 2.820 1430.070 2.960 ;
        RECT 1428.370 2.760 1428.690 2.820 ;
        RECT 1429.750 2.760 1430.070 2.820 ;
      LAYER via ;
        RECT 1291.320 1655.840 1291.580 1656.100 ;
        RECT 1296.840 1655.840 1297.100 1656.100 ;
        RECT 1291.320 1577.300 1291.580 1577.560 ;
        RECT 1428.400 1577.300 1428.660 1577.560 ;
        RECT 1428.400 2.760 1428.660 3.020 ;
        RECT 1429.780 2.760 1430.040 3.020 ;
      LAYER met2 ;
        RECT 1296.740 1700.340 1297.020 1704.000 ;
        RECT 1296.740 1700.000 1297.040 1700.340 ;
        RECT 1296.900 1656.130 1297.040 1700.000 ;
        RECT 1291.320 1655.810 1291.580 1656.130 ;
        RECT 1296.840 1655.810 1297.100 1656.130 ;
        RECT 1291.380 1577.590 1291.520 1655.810 ;
        RECT 1291.320 1577.270 1291.580 1577.590 ;
        RECT 1428.400 1577.270 1428.660 1577.590 ;
        RECT 1428.460 3.050 1428.600 1577.270 ;
        RECT 1428.400 2.730 1428.660 3.050 ;
        RECT 1429.780 2.730 1430.040 3.050 ;
        RECT 1429.840 2.400 1429.980 2.730 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1366.345 1685.465 1366.515 1689.715 ;
        RECT 1404.065 1687.845 1404.235 1689.715 ;
      LAYER mcon ;
        RECT 1366.345 1689.545 1366.515 1689.715 ;
        RECT 1404.065 1689.545 1404.235 1689.715 ;
      LAYER met1 ;
        RECT 1366.285 1689.700 1366.575 1689.745 ;
        RECT 1404.005 1689.700 1404.295 1689.745 ;
        RECT 1366.285 1689.560 1404.295 1689.700 ;
        RECT 1366.285 1689.515 1366.575 1689.560 ;
        RECT 1404.005 1689.515 1404.295 1689.560 ;
        RECT 1403.990 1688.000 1404.310 1688.060 ;
        RECT 1403.795 1687.860 1404.310 1688.000 ;
        RECT 1403.990 1687.800 1404.310 1687.860 ;
        RECT 1298.650 1685.620 1298.970 1685.680 ;
        RECT 1318.430 1685.620 1318.750 1685.680 ;
        RECT 1298.650 1685.480 1318.750 1685.620 ;
        RECT 1298.650 1685.420 1298.970 1685.480 ;
        RECT 1318.430 1685.420 1318.750 1685.480 ;
        RECT 1338.670 1685.620 1338.990 1685.680 ;
        RECT 1366.285 1685.620 1366.575 1685.665 ;
        RECT 1338.670 1685.480 1366.575 1685.620 ;
        RECT 1338.670 1685.420 1338.990 1685.480 ;
        RECT 1366.285 1685.435 1366.575 1685.480 ;
        RECT 1403.990 1678.280 1404.310 1678.540 ;
        RECT 1404.080 1678.140 1404.220 1678.280 ;
        RECT 1403.620 1678.000 1404.220 1678.140 ;
        RECT 1403.620 1677.520 1403.760 1678.000 ;
        RECT 1403.530 1677.260 1403.850 1677.520 ;
        RECT 1403.990 34.580 1404.310 34.640 ;
        RECT 1447.690 34.580 1448.010 34.640 ;
        RECT 1403.990 34.440 1448.010 34.580 ;
        RECT 1403.990 34.380 1404.310 34.440 ;
        RECT 1447.690 34.380 1448.010 34.440 ;
      LAYER via ;
        RECT 1404.020 1687.800 1404.280 1688.060 ;
        RECT 1298.680 1685.420 1298.940 1685.680 ;
        RECT 1318.460 1685.420 1318.720 1685.680 ;
        RECT 1338.700 1685.420 1338.960 1685.680 ;
        RECT 1404.020 1678.280 1404.280 1678.540 ;
        RECT 1403.560 1677.260 1403.820 1677.520 ;
        RECT 1404.020 34.380 1404.280 34.640 ;
        RECT 1447.720 34.380 1447.980 34.640 ;
      LAYER met2 ;
        RECT 1298.580 1700.340 1298.860 1704.000 ;
        RECT 1298.580 1700.000 1298.880 1700.340 ;
        RECT 1298.740 1685.710 1298.880 1700.000 ;
        RECT 1404.020 1687.770 1404.280 1688.090 ;
        RECT 1298.680 1685.390 1298.940 1685.710 ;
        RECT 1318.460 1685.565 1318.720 1685.710 ;
        RECT 1338.700 1685.565 1338.960 1685.710 ;
        RECT 1318.450 1685.195 1318.730 1685.565 ;
        RECT 1338.690 1685.195 1338.970 1685.565 ;
        RECT 1404.080 1678.570 1404.220 1687.770 ;
        RECT 1404.020 1678.250 1404.280 1678.570 ;
        RECT 1403.560 1677.230 1403.820 1677.550 ;
        RECT 1403.620 1631.730 1403.760 1677.230 ;
        RECT 1403.620 1631.590 1404.220 1631.730 ;
        RECT 1404.080 34.670 1404.220 1631.590 ;
        RECT 1404.020 34.350 1404.280 34.670 ;
        RECT 1447.720 34.350 1447.980 34.670 ;
        RECT 1447.780 2.400 1447.920 34.350 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
      LAYER via2 ;
        RECT 1318.450 1685.240 1318.730 1685.520 ;
        RECT 1338.690 1685.240 1338.970 1685.520 ;
      LAYER met3 ;
        RECT 1318.425 1685.530 1318.755 1685.545 ;
        RECT 1338.665 1685.530 1338.995 1685.545 ;
        RECT 1318.425 1685.230 1338.995 1685.530 ;
        RECT 1318.425 1685.215 1318.755 1685.230 ;
        RECT 1338.665 1685.215 1338.995 1685.230 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1300.490 1685.960 1300.810 1686.020 ;
        RECT 1303.710 1685.960 1304.030 1686.020 ;
        RECT 1300.490 1685.820 1304.030 1685.960 ;
        RECT 1300.490 1685.760 1300.810 1685.820 ;
        RECT 1303.710 1685.760 1304.030 1685.820 ;
        RECT 1303.710 1675.420 1304.030 1675.480 ;
        RECT 1462.870 1675.420 1463.190 1675.480 ;
        RECT 1303.710 1675.280 1463.190 1675.420 ;
        RECT 1303.710 1675.220 1304.030 1675.280 ;
        RECT 1462.870 1675.220 1463.190 1675.280 ;
      LAYER via ;
        RECT 1300.520 1685.760 1300.780 1686.020 ;
        RECT 1303.740 1685.760 1304.000 1686.020 ;
        RECT 1303.740 1675.220 1304.000 1675.480 ;
        RECT 1462.900 1675.220 1463.160 1675.480 ;
      LAYER met2 ;
        RECT 1300.420 1700.340 1300.700 1704.000 ;
        RECT 1300.420 1700.000 1300.720 1700.340 ;
        RECT 1300.580 1686.050 1300.720 1700.000 ;
        RECT 1300.520 1685.730 1300.780 1686.050 ;
        RECT 1303.740 1685.730 1304.000 1686.050 ;
        RECT 1303.800 1675.510 1303.940 1685.730 ;
        RECT 1303.740 1675.190 1304.000 1675.510 ;
        RECT 1462.900 1675.190 1463.160 1675.510 ;
        RECT 1462.960 17.410 1463.100 1675.190 ;
        RECT 1462.960 17.270 1465.860 17.410 ;
        RECT 1465.720 2.400 1465.860 17.270 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1302.330 1661.820 1302.650 1661.880 ;
        RECT 1484.030 1661.820 1484.350 1661.880 ;
        RECT 1302.330 1661.680 1484.350 1661.820 ;
        RECT 1302.330 1661.620 1302.650 1661.680 ;
        RECT 1484.030 1661.620 1484.350 1661.680 ;
      LAYER via ;
        RECT 1302.360 1661.620 1302.620 1661.880 ;
        RECT 1484.060 1661.620 1484.320 1661.880 ;
      LAYER met2 ;
        RECT 1302.260 1700.340 1302.540 1704.000 ;
        RECT 1302.260 1700.000 1302.560 1700.340 ;
        RECT 1302.420 1661.910 1302.560 1700.000 ;
        RECT 1302.360 1661.590 1302.620 1661.910 ;
        RECT 1484.060 1661.590 1484.320 1661.910 ;
        RECT 1484.120 7.210 1484.260 1661.590 ;
        RECT 1483.660 7.070 1484.260 7.210 ;
        RECT 1483.660 2.400 1483.800 7.070 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1304.630 1640.740 1304.950 1640.800 ;
        RECT 1497.370 1640.740 1497.690 1640.800 ;
        RECT 1304.630 1640.600 1497.690 1640.740 ;
        RECT 1304.630 1640.540 1304.950 1640.600 ;
        RECT 1497.370 1640.540 1497.690 1640.600 ;
        RECT 1497.370 2.960 1497.690 3.020 ;
        RECT 1501.510 2.960 1501.830 3.020 ;
        RECT 1497.370 2.820 1501.830 2.960 ;
        RECT 1497.370 2.760 1497.690 2.820 ;
        RECT 1501.510 2.760 1501.830 2.820 ;
      LAYER via ;
        RECT 1304.660 1640.540 1304.920 1640.800 ;
        RECT 1497.400 1640.540 1497.660 1640.800 ;
        RECT 1497.400 2.760 1497.660 3.020 ;
        RECT 1501.540 2.760 1501.800 3.020 ;
      LAYER met2 ;
        RECT 1304.100 1700.340 1304.380 1704.000 ;
        RECT 1304.100 1700.000 1304.400 1700.340 ;
        RECT 1304.260 1667.770 1304.400 1700.000 ;
        RECT 1303.800 1667.630 1304.400 1667.770 ;
        RECT 1303.800 1666.410 1303.940 1667.630 ;
        RECT 1303.800 1666.270 1304.860 1666.410 ;
        RECT 1304.720 1640.830 1304.860 1666.270 ;
        RECT 1304.660 1640.510 1304.920 1640.830 ;
        RECT 1497.400 1640.510 1497.660 1640.830 ;
        RECT 1497.460 3.050 1497.600 1640.510 ;
        RECT 1497.400 2.730 1497.660 3.050 ;
        RECT 1501.540 2.730 1501.800 3.050 ;
        RECT 1501.600 2.400 1501.740 2.730 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1306.010 1684.600 1306.330 1684.660 ;
        RECT 1309.230 1684.600 1309.550 1684.660 ;
        RECT 1306.010 1684.460 1309.550 1684.600 ;
        RECT 1306.010 1684.400 1306.330 1684.460 ;
        RECT 1309.230 1684.400 1309.550 1684.460 ;
        RECT 1309.230 1626.460 1309.550 1626.520 ;
        RECT 1518.070 1626.460 1518.390 1626.520 ;
        RECT 1309.230 1626.320 1518.390 1626.460 ;
        RECT 1309.230 1626.260 1309.550 1626.320 ;
        RECT 1518.070 1626.260 1518.390 1626.320 ;
        RECT 1518.070 2.960 1518.390 3.020 ;
        RECT 1518.990 2.960 1519.310 3.020 ;
        RECT 1518.070 2.820 1519.310 2.960 ;
        RECT 1518.070 2.760 1518.390 2.820 ;
        RECT 1518.990 2.760 1519.310 2.820 ;
      LAYER via ;
        RECT 1306.040 1684.400 1306.300 1684.660 ;
        RECT 1309.260 1684.400 1309.520 1684.660 ;
        RECT 1309.260 1626.260 1309.520 1626.520 ;
        RECT 1518.100 1626.260 1518.360 1626.520 ;
        RECT 1518.100 2.760 1518.360 3.020 ;
        RECT 1519.020 2.760 1519.280 3.020 ;
      LAYER met2 ;
        RECT 1305.940 1700.340 1306.220 1704.000 ;
        RECT 1305.940 1700.000 1306.240 1700.340 ;
        RECT 1306.100 1684.690 1306.240 1700.000 ;
        RECT 1306.040 1684.370 1306.300 1684.690 ;
        RECT 1309.260 1684.370 1309.520 1684.690 ;
        RECT 1309.320 1626.550 1309.460 1684.370 ;
        RECT 1309.260 1626.230 1309.520 1626.550 ;
        RECT 1518.100 1626.230 1518.360 1626.550 ;
        RECT 1518.160 3.050 1518.300 1626.230 ;
        RECT 1518.100 2.730 1518.360 3.050 ;
        RECT 1519.020 2.730 1519.280 3.050 ;
        RECT 1519.080 2.400 1519.220 2.730 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 717.210 1576.820 717.530 1576.880 ;
        RECT 1224.130 1576.820 1224.450 1576.880 ;
        RECT 717.210 1576.680 1224.450 1576.820 ;
        RECT 717.210 1576.620 717.530 1576.680 ;
        RECT 1224.130 1576.620 1224.450 1576.680 ;
      LAYER via ;
        RECT 717.240 1576.620 717.500 1576.880 ;
        RECT 1224.160 1576.620 1224.420 1576.880 ;
      LAYER met2 ;
        RECT 1223.140 1700.410 1223.420 1704.000 ;
        RECT 1223.140 1700.270 1223.900 1700.410 ;
        RECT 1223.140 1700.000 1223.420 1700.270 ;
        RECT 1223.760 1677.970 1223.900 1700.270 ;
        RECT 1223.760 1677.830 1224.360 1677.970 ;
        RECT 1224.220 1576.910 1224.360 1677.830 ;
        RECT 717.240 1576.590 717.500 1576.910 ;
        RECT 1224.160 1576.590 1224.420 1576.910 ;
        RECT 717.300 16.730 717.440 1576.590 ;
        RECT 716.380 16.590 717.440 16.730 ;
        RECT 716.380 2.400 716.520 16.590 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1308.310 1631.360 1308.630 1631.620 ;
        RECT 1308.400 1630.600 1308.540 1631.360 ;
        RECT 1308.310 1630.340 1308.630 1630.600 ;
        RECT 1308.310 1598.580 1308.630 1598.640 ;
        RECT 1531.870 1598.580 1532.190 1598.640 ;
        RECT 1308.310 1598.440 1532.190 1598.580 ;
        RECT 1308.310 1598.380 1308.630 1598.440 ;
        RECT 1531.870 1598.380 1532.190 1598.440 ;
      LAYER via ;
        RECT 1308.340 1631.360 1308.600 1631.620 ;
        RECT 1308.340 1630.340 1308.600 1630.600 ;
        RECT 1308.340 1598.380 1308.600 1598.640 ;
        RECT 1531.900 1598.380 1532.160 1598.640 ;
      LAYER met2 ;
        RECT 1307.780 1700.340 1308.060 1704.000 ;
        RECT 1307.780 1700.000 1308.080 1700.340 ;
        RECT 1307.940 1668.450 1308.080 1700.000 ;
        RECT 1307.940 1668.310 1308.540 1668.450 ;
        RECT 1308.400 1631.650 1308.540 1668.310 ;
        RECT 1308.340 1631.330 1308.600 1631.650 ;
        RECT 1308.340 1630.310 1308.600 1630.630 ;
        RECT 1308.400 1598.670 1308.540 1630.310 ;
        RECT 1308.340 1598.350 1308.600 1598.670 ;
        RECT 1531.900 1598.350 1532.160 1598.670 ;
        RECT 1531.960 17.410 1532.100 1598.350 ;
        RECT 1531.960 17.270 1537.160 17.410 ;
        RECT 1537.020 2.400 1537.160 17.270 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1309.690 1656.380 1310.010 1656.440 ;
        RECT 1304.260 1656.240 1310.010 1656.380 ;
        RECT 1304.260 1656.100 1304.400 1656.240 ;
        RECT 1309.690 1656.180 1310.010 1656.240 ;
        RECT 1304.170 1655.840 1304.490 1656.100 ;
        RECT 1304.170 1556.760 1304.490 1556.820 ;
        RECT 1552.570 1556.760 1552.890 1556.820 ;
        RECT 1304.170 1556.620 1552.890 1556.760 ;
        RECT 1304.170 1556.560 1304.490 1556.620 ;
        RECT 1552.570 1556.560 1552.890 1556.620 ;
      LAYER via ;
        RECT 1309.720 1656.180 1309.980 1656.440 ;
        RECT 1304.200 1655.840 1304.460 1656.100 ;
        RECT 1304.200 1556.560 1304.460 1556.820 ;
        RECT 1552.600 1556.560 1552.860 1556.820 ;
      LAYER met2 ;
        RECT 1309.620 1700.340 1309.900 1704.000 ;
        RECT 1309.620 1700.000 1309.920 1700.340 ;
        RECT 1309.780 1656.470 1309.920 1700.000 ;
        RECT 1309.720 1656.150 1309.980 1656.470 ;
        RECT 1304.200 1655.810 1304.460 1656.130 ;
        RECT 1304.260 1556.850 1304.400 1655.810 ;
        RECT 1304.200 1556.530 1304.460 1556.850 ;
        RECT 1552.600 1556.530 1552.860 1556.850 ;
        RECT 1552.660 17.410 1552.800 1556.530 ;
        RECT 1552.660 17.270 1555.100 17.410 ;
        RECT 1554.960 2.400 1555.100 17.270 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1311.530 1619.660 1311.850 1619.720 ;
        RECT 1566.830 1619.660 1567.150 1619.720 ;
        RECT 1311.530 1619.520 1567.150 1619.660 ;
        RECT 1311.530 1619.460 1311.850 1619.520 ;
        RECT 1566.830 1619.460 1567.150 1619.520 ;
        RECT 1566.830 20.980 1567.150 21.040 ;
        RECT 1572.810 20.980 1573.130 21.040 ;
        RECT 1566.830 20.840 1573.130 20.980 ;
        RECT 1566.830 20.780 1567.150 20.840 ;
        RECT 1572.810 20.780 1573.130 20.840 ;
      LAYER via ;
        RECT 1311.560 1619.460 1311.820 1619.720 ;
        RECT 1566.860 1619.460 1567.120 1619.720 ;
        RECT 1566.860 20.780 1567.120 21.040 ;
        RECT 1572.840 20.780 1573.100 21.040 ;
      LAYER met2 ;
        RECT 1311.460 1700.340 1311.740 1704.000 ;
        RECT 1311.460 1700.000 1311.760 1700.340 ;
        RECT 1311.620 1619.750 1311.760 1700.000 ;
        RECT 1311.560 1619.430 1311.820 1619.750 ;
        RECT 1566.860 1619.430 1567.120 1619.750 ;
        RECT 1566.920 21.070 1567.060 1619.430 ;
        RECT 1566.860 20.750 1567.120 21.070 ;
        RECT 1572.840 20.750 1573.100 21.070 ;
        RECT 1572.900 2.400 1573.040 20.750 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1313.370 1656.720 1313.690 1656.780 ;
        RECT 1313.370 1656.580 1316.360 1656.720 ;
        RECT 1313.370 1656.520 1313.690 1656.580 ;
        RECT 1316.220 1656.440 1316.360 1656.580 ;
        RECT 1316.130 1656.180 1316.450 1656.440 ;
        RECT 1316.130 1549.960 1316.450 1550.020 ;
        RECT 1587.070 1549.960 1587.390 1550.020 ;
        RECT 1316.130 1549.820 1587.390 1549.960 ;
        RECT 1316.130 1549.760 1316.450 1549.820 ;
        RECT 1587.070 1549.760 1587.390 1549.820 ;
      LAYER via ;
        RECT 1313.400 1656.520 1313.660 1656.780 ;
        RECT 1316.160 1656.180 1316.420 1656.440 ;
        RECT 1316.160 1549.760 1316.420 1550.020 ;
        RECT 1587.100 1549.760 1587.360 1550.020 ;
      LAYER met2 ;
        RECT 1313.300 1700.340 1313.580 1704.000 ;
        RECT 1313.300 1700.000 1313.600 1700.340 ;
        RECT 1313.460 1656.810 1313.600 1700.000 ;
        RECT 1313.400 1656.490 1313.660 1656.810 ;
        RECT 1316.160 1656.150 1316.420 1656.470 ;
        RECT 1316.220 1550.050 1316.360 1656.150 ;
        RECT 1316.160 1549.730 1316.420 1550.050 ;
        RECT 1587.100 1549.730 1587.360 1550.050 ;
        RECT 1587.160 17.410 1587.300 1549.730 ;
        RECT 1587.160 17.270 1590.520 17.410 ;
        RECT 1590.380 2.400 1590.520 17.270 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1315.210 1612.180 1315.530 1612.240 ;
        RECT 1607.770 1612.180 1608.090 1612.240 ;
        RECT 1315.210 1612.040 1608.090 1612.180 ;
        RECT 1315.210 1611.980 1315.530 1612.040 ;
        RECT 1607.770 1611.980 1608.090 1612.040 ;
      LAYER via ;
        RECT 1315.240 1611.980 1315.500 1612.240 ;
        RECT 1607.800 1611.980 1608.060 1612.240 ;
      LAYER met2 ;
        RECT 1315.140 1700.340 1315.420 1704.000 ;
        RECT 1315.140 1700.000 1315.440 1700.340 ;
        RECT 1315.300 1612.270 1315.440 1700.000 ;
        RECT 1315.240 1611.950 1315.500 1612.270 ;
        RECT 1607.800 1611.950 1608.060 1612.270 ;
        RECT 1607.860 17.410 1608.000 1611.950 ;
        RECT 1607.860 17.270 1608.460 17.410 ;
        RECT 1608.320 2.400 1608.460 17.270 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1312.910 1678.820 1313.230 1678.880 ;
        RECT 1317.050 1678.820 1317.370 1678.880 ;
        RECT 1312.910 1678.680 1317.370 1678.820 ;
        RECT 1312.910 1678.620 1313.230 1678.680 ;
        RECT 1317.050 1678.620 1317.370 1678.680 ;
        RECT 1312.450 1466.660 1312.770 1466.720 ;
        RECT 1621.570 1466.660 1621.890 1466.720 ;
        RECT 1312.450 1466.520 1621.890 1466.660 ;
        RECT 1312.450 1466.460 1312.770 1466.520 ;
        RECT 1621.570 1466.460 1621.890 1466.520 ;
      LAYER via ;
        RECT 1312.940 1678.620 1313.200 1678.880 ;
        RECT 1317.080 1678.620 1317.340 1678.880 ;
        RECT 1312.480 1466.460 1312.740 1466.720 ;
        RECT 1621.600 1466.460 1621.860 1466.720 ;
      LAYER met2 ;
        RECT 1316.980 1700.340 1317.260 1704.000 ;
        RECT 1316.980 1700.000 1317.280 1700.340 ;
        RECT 1317.140 1678.910 1317.280 1700.000 ;
        RECT 1312.940 1678.590 1313.200 1678.910 ;
        RECT 1317.080 1678.590 1317.340 1678.910 ;
        RECT 1313.000 1659.610 1313.140 1678.590 ;
        RECT 1312.540 1659.470 1313.140 1659.610 ;
        RECT 1312.540 1466.750 1312.680 1659.470 ;
        RECT 1312.480 1466.430 1312.740 1466.750 ;
        RECT 1621.600 1466.430 1621.860 1466.750 ;
        RECT 1621.660 17.410 1621.800 1466.430 ;
        RECT 1621.660 17.270 1626.400 17.410 ;
        RECT 1626.260 2.400 1626.400 17.270 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1318.890 1684.940 1319.210 1685.000 ;
        RECT 1322.110 1684.940 1322.430 1685.000 ;
        RECT 1318.890 1684.800 1322.430 1684.940 ;
        RECT 1318.890 1684.740 1319.210 1684.800 ;
        RECT 1322.110 1684.740 1322.430 1684.800 ;
        RECT 1322.110 1640.400 1322.430 1640.460 ;
        RECT 1642.270 1640.400 1642.590 1640.460 ;
        RECT 1322.110 1640.260 1642.590 1640.400 ;
        RECT 1322.110 1640.200 1322.430 1640.260 ;
        RECT 1642.270 1640.200 1642.590 1640.260 ;
        RECT 1642.270 1140.400 1642.590 1140.660 ;
        RECT 1642.360 1139.640 1642.500 1140.400 ;
        RECT 1642.270 1139.380 1642.590 1139.640 ;
        RECT 1642.270 381.520 1642.590 381.780 ;
        RECT 1642.360 380.760 1642.500 381.520 ;
        RECT 1642.270 380.500 1642.590 380.760 ;
      LAYER via ;
        RECT 1318.920 1684.740 1319.180 1685.000 ;
        RECT 1322.140 1684.740 1322.400 1685.000 ;
        RECT 1322.140 1640.200 1322.400 1640.460 ;
        RECT 1642.300 1640.200 1642.560 1640.460 ;
        RECT 1642.300 1140.400 1642.560 1140.660 ;
        RECT 1642.300 1139.380 1642.560 1139.640 ;
        RECT 1642.300 381.520 1642.560 381.780 ;
        RECT 1642.300 380.500 1642.560 380.760 ;
      LAYER met2 ;
        RECT 1318.820 1700.340 1319.100 1704.000 ;
        RECT 1318.820 1700.000 1319.120 1700.340 ;
        RECT 1318.980 1685.030 1319.120 1700.000 ;
        RECT 1318.920 1684.710 1319.180 1685.030 ;
        RECT 1322.140 1684.710 1322.400 1685.030 ;
        RECT 1322.200 1640.490 1322.340 1684.710 ;
        RECT 1322.140 1640.170 1322.400 1640.490 ;
        RECT 1642.300 1640.170 1642.560 1640.490 ;
        RECT 1642.360 1140.690 1642.500 1640.170 ;
        RECT 1642.300 1140.370 1642.560 1140.690 ;
        RECT 1642.300 1139.350 1642.560 1139.670 ;
        RECT 1642.360 381.810 1642.500 1139.350 ;
        RECT 1642.300 381.490 1642.560 381.810 ;
        RECT 1642.300 380.470 1642.560 380.790 ;
        RECT 1642.360 17.410 1642.500 380.470 ;
        RECT 1642.360 17.270 1644.340 17.410 ;
        RECT 1644.200 2.400 1644.340 17.270 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1412.805 1684.105 1412.975 1688.355 ;
      LAYER mcon ;
        RECT 1412.805 1688.185 1412.975 1688.355 ;
      LAYER met1 ;
        RECT 1320.730 1689.020 1321.050 1689.080 ;
        RECT 1320.730 1688.880 1363.280 1689.020 ;
        RECT 1320.730 1688.820 1321.050 1688.880 ;
        RECT 1363.140 1688.340 1363.280 1688.880 ;
        RECT 1412.745 1688.340 1413.035 1688.385 ;
        RECT 1363.140 1688.200 1413.035 1688.340 ;
        RECT 1412.745 1688.155 1413.035 1688.200 ;
        RECT 1414.570 1685.960 1414.890 1686.020 ;
        RECT 1416.410 1685.960 1416.730 1686.020 ;
        RECT 1414.570 1685.820 1416.730 1685.960 ;
        RECT 1414.570 1685.760 1414.890 1685.820 ;
        RECT 1416.410 1685.760 1416.730 1685.820 ;
        RECT 1412.745 1684.260 1413.035 1684.305 ;
        RECT 1414.570 1684.260 1414.890 1684.320 ;
        RECT 1412.745 1684.120 1414.890 1684.260 ;
        RECT 1412.745 1684.075 1413.035 1684.120 ;
        RECT 1414.570 1684.060 1414.890 1684.120 ;
        RECT 1417.790 24.720 1418.110 24.780 ;
        RECT 1417.790 24.580 1459.420 24.720 ;
        RECT 1417.790 24.520 1418.110 24.580 ;
        RECT 1459.280 24.380 1459.420 24.580 ;
        RECT 1662.050 24.380 1662.370 24.440 ;
        RECT 1459.280 24.240 1662.370 24.380 ;
        RECT 1662.050 24.180 1662.370 24.240 ;
      LAYER via ;
        RECT 1320.760 1688.820 1321.020 1689.080 ;
        RECT 1414.600 1685.760 1414.860 1686.020 ;
        RECT 1416.440 1685.760 1416.700 1686.020 ;
        RECT 1414.600 1684.060 1414.860 1684.320 ;
        RECT 1417.820 24.520 1418.080 24.780 ;
        RECT 1662.080 24.180 1662.340 24.440 ;
      LAYER met2 ;
        RECT 1320.660 1700.340 1320.940 1704.000 ;
        RECT 1320.660 1700.000 1320.960 1700.340 ;
        RECT 1320.820 1689.110 1320.960 1700.000 ;
        RECT 1320.760 1688.790 1321.020 1689.110 ;
        RECT 1414.600 1685.730 1414.860 1686.050 ;
        RECT 1416.440 1685.730 1416.700 1686.050 ;
        RECT 1414.660 1684.350 1414.800 1685.730 ;
        RECT 1416.500 1685.450 1416.640 1685.730 ;
        RECT 1416.500 1685.310 1417.100 1685.450 ;
        RECT 1414.600 1684.030 1414.860 1684.350 ;
        RECT 1416.960 1676.610 1417.100 1685.310 ;
        RECT 1416.960 1676.470 1418.020 1676.610 ;
        RECT 1417.880 24.810 1418.020 1676.470 ;
        RECT 1417.820 24.490 1418.080 24.810 ;
        RECT 1662.080 24.150 1662.340 24.470 ;
        RECT 1662.140 2.400 1662.280 24.150 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1322.570 1591.440 1322.890 1591.500 ;
        RECT 1676.770 1591.440 1677.090 1591.500 ;
        RECT 1322.570 1591.300 1677.090 1591.440 ;
        RECT 1322.570 1591.240 1322.890 1591.300 ;
        RECT 1676.770 1591.240 1677.090 1591.300 ;
      LAYER via ;
        RECT 1322.600 1591.240 1322.860 1591.500 ;
        RECT 1676.800 1591.240 1677.060 1591.500 ;
      LAYER met2 ;
        RECT 1322.500 1700.340 1322.780 1704.000 ;
        RECT 1322.500 1700.000 1322.800 1700.340 ;
        RECT 1322.660 1591.530 1322.800 1700.000 ;
        RECT 1322.600 1591.210 1322.860 1591.530 ;
        RECT 1676.800 1591.210 1677.060 1591.530 ;
        RECT 1676.860 17.410 1677.000 1591.210 ;
        RECT 1676.860 17.270 1679.760 17.410 ;
        RECT 1679.620 2.400 1679.760 17.270 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1319.810 1685.620 1320.130 1685.680 ;
        RECT 1324.410 1685.620 1324.730 1685.680 ;
        RECT 1319.810 1685.480 1324.730 1685.620 ;
        RECT 1319.810 1685.420 1320.130 1685.480 ;
        RECT 1324.410 1685.420 1324.730 1685.480 ;
        RECT 1319.810 1542.820 1320.130 1542.880 ;
        RECT 1697.470 1542.820 1697.790 1542.880 ;
        RECT 1319.810 1542.680 1697.790 1542.820 ;
        RECT 1319.810 1542.620 1320.130 1542.680 ;
        RECT 1697.470 1542.620 1697.790 1542.680 ;
      LAYER via ;
        RECT 1319.840 1685.420 1320.100 1685.680 ;
        RECT 1324.440 1685.420 1324.700 1685.680 ;
        RECT 1319.840 1542.620 1320.100 1542.880 ;
        RECT 1697.500 1542.620 1697.760 1542.880 ;
      LAYER met2 ;
        RECT 1324.340 1700.340 1324.620 1704.000 ;
        RECT 1324.340 1700.000 1324.640 1700.340 ;
        RECT 1324.500 1685.710 1324.640 1700.000 ;
        RECT 1319.840 1685.390 1320.100 1685.710 ;
        RECT 1324.440 1685.390 1324.700 1685.710 ;
        RECT 1319.900 1542.910 1320.040 1685.390 ;
        RECT 1319.840 1542.590 1320.100 1542.910 ;
        RECT 1697.500 1542.590 1697.760 1542.910 ;
        RECT 1697.560 2.400 1697.700 1542.590 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 737.910 1570.020 738.230 1570.080 ;
        RECT 1225.050 1570.020 1225.370 1570.080 ;
        RECT 737.910 1569.880 1225.370 1570.020 ;
        RECT 737.910 1569.820 738.230 1569.880 ;
        RECT 1225.050 1569.820 1225.370 1569.880 ;
      LAYER via ;
        RECT 737.940 1569.820 738.200 1570.080 ;
        RECT 1225.080 1569.820 1225.340 1570.080 ;
      LAYER met2 ;
        RECT 1224.980 1700.340 1225.260 1704.000 ;
        RECT 1224.980 1700.000 1225.280 1700.340 ;
        RECT 1225.140 1570.110 1225.280 1700.000 ;
        RECT 737.940 1569.790 738.200 1570.110 ;
        RECT 1225.080 1569.790 1225.340 1570.110 ;
        RECT 738.000 16.730 738.140 1569.790 ;
        RECT 734.320 16.590 738.140 16.730 ;
        RECT 734.320 2.400 734.460 16.590 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1328.165 1683.765 1328.335 1688.695 ;
      LAYER mcon ;
        RECT 1328.165 1688.525 1328.335 1688.695 ;
      LAYER met1 ;
        RECT 1326.250 1688.680 1326.570 1688.740 ;
        RECT 1328.105 1688.680 1328.395 1688.725 ;
        RECT 1326.250 1688.540 1328.395 1688.680 ;
        RECT 1326.250 1688.480 1326.570 1688.540 ;
        RECT 1328.105 1688.495 1328.395 1688.540 ;
        RECT 1328.090 1683.920 1328.410 1683.980 ;
        RECT 1328.090 1683.780 1328.605 1683.920 ;
        RECT 1328.090 1683.720 1328.410 1683.780 ;
        RECT 1328.090 1646.860 1328.410 1646.920 ;
        RECT 1711.270 1646.860 1711.590 1646.920 ;
        RECT 1328.090 1646.720 1711.590 1646.860 ;
        RECT 1328.090 1646.660 1328.410 1646.720 ;
        RECT 1711.270 1646.660 1711.590 1646.720 ;
      LAYER via ;
        RECT 1326.280 1688.480 1326.540 1688.740 ;
        RECT 1328.120 1683.720 1328.380 1683.980 ;
        RECT 1328.120 1646.660 1328.380 1646.920 ;
        RECT 1711.300 1646.660 1711.560 1646.920 ;
      LAYER met2 ;
        RECT 1326.180 1700.340 1326.460 1704.000 ;
        RECT 1326.180 1700.000 1326.480 1700.340 ;
        RECT 1326.340 1688.770 1326.480 1700.000 ;
        RECT 1326.280 1688.450 1326.540 1688.770 ;
        RECT 1328.120 1683.690 1328.380 1684.010 ;
        RECT 1328.180 1646.950 1328.320 1683.690 ;
        RECT 1328.120 1646.630 1328.380 1646.950 ;
        RECT 1711.300 1646.630 1711.560 1646.950 ;
        RECT 1711.360 17.410 1711.500 1646.630 ;
        RECT 1711.360 17.270 1715.640 17.410 ;
        RECT 1715.500 2.400 1715.640 17.270 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1449.605 1687.165 1450.695 1687.335 ;
      LAYER mcon ;
        RECT 1450.525 1687.165 1450.695 1687.335 ;
      LAYER met1 ;
        RECT 1328.090 1687.320 1328.410 1687.380 ;
        RECT 1449.545 1687.320 1449.835 1687.365 ;
        RECT 1328.090 1687.180 1449.835 1687.320 ;
        RECT 1328.090 1687.120 1328.410 1687.180 ;
        RECT 1449.545 1687.135 1449.835 1687.180 ;
        RECT 1450.465 1687.320 1450.755 1687.365 ;
        RECT 1731.970 1687.320 1732.290 1687.380 ;
        RECT 1450.465 1687.180 1732.290 1687.320 ;
        RECT 1450.465 1687.135 1450.755 1687.180 ;
        RECT 1731.970 1687.120 1732.290 1687.180 ;
      LAYER via ;
        RECT 1328.120 1687.120 1328.380 1687.380 ;
        RECT 1732.000 1687.120 1732.260 1687.380 ;
      LAYER met2 ;
        RECT 1328.020 1700.340 1328.300 1704.000 ;
        RECT 1328.020 1700.000 1328.320 1700.340 ;
        RECT 1328.180 1687.410 1328.320 1700.000 ;
        RECT 1328.120 1687.090 1328.380 1687.410 ;
        RECT 1732.000 1687.090 1732.260 1687.410 ;
        RECT 1732.060 17.410 1732.200 1687.090 ;
        RECT 1732.060 17.270 1733.580 17.410 ;
        RECT 1733.440 2.400 1733.580 17.270 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1329.930 1681.540 1330.250 1681.600 ;
        RECT 1745.770 1681.540 1746.090 1681.600 ;
        RECT 1329.930 1681.400 1746.090 1681.540 ;
        RECT 1329.930 1681.340 1330.250 1681.400 ;
        RECT 1745.770 1681.340 1746.090 1681.400 ;
      LAYER via ;
        RECT 1329.960 1681.340 1330.220 1681.600 ;
        RECT 1745.800 1681.340 1746.060 1681.600 ;
      LAYER met2 ;
        RECT 1329.860 1700.340 1330.140 1704.000 ;
        RECT 1329.860 1700.000 1330.160 1700.340 ;
        RECT 1330.020 1681.630 1330.160 1700.000 ;
        RECT 1329.960 1681.310 1330.220 1681.630 ;
        RECT 1745.800 1681.310 1746.060 1681.630 ;
        RECT 1745.860 17.410 1746.000 1681.310 ;
        RECT 1745.860 17.270 1751.520 17.410 ;
        RECT 1751.380 2.400 1751.520 17.270 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1334.145 1674.245 1334.315 1683.595 ;
      LAYER mcon ;
        RECT 1334.145 1683.425 1334.315 1683.595 ;
      LAYER met1 ;
        RECT 1331.770 1687.660 1332.090 1687.720 ;
        RECT 1333.150 1687.660 1333.470 1687.720 ;
        RECT 1331.770 1687.520 1333.470 1687.660 ;
        RECT 1331.770 1687.460 1332.090 1687.520 ;
        RECT 1333.150 1687.460 1333.470 1687.520 ;
        RECT 1333.150 1683.920 1333.470 1683.980 ;
        RECT 1333.150 1683.780 1334.300 1683.920 ;
        RECT 1333.150 1683.720 1333.470 1683.780 ;
        RECT 1334.160 1683.625 1334.300 1683.780 ;
        RECT 1334.085 1683.580 1334.375 1683.625 ;
        RECT 1334.085 1683.440 1334.485 1683.580 ;
        RECT 1334.085 1683.395 1334.375 1683.440 ;
        RECT 1334.085 1674.400 1334.375 1674.445 ;
        RECT 1766.470 1674.400 1766.790 1674.460 ;
        RECT 1334.085 1674.260 1766.790 1674.400 ;
        RECT 1334.085 1674.215 1334.375 1674.260 ;
        RECT 1766.470 1674.200 1766.790 1674.260 ;
      LAYER via ;
        RECT 1331.800 1687.460 1332.060 1687.720 ;
        RECT 1333.180 1687.460 1333.440 1687.720 ;
        RECT 1333.180 1683.720 1333.440 1683.980 ;
        RECT 1766.500 1674.200 1766.760 1674.460 ;
      LAYER met2 ;
        RECT 1331.700 1700.340 1331.980 1704.000 ;
        RECT 1331.700 1700.000 1332.000 1700.340 ;
        RECT 1331.860 1687.750 1332.000 1700.000 ;
        RECT 1331.800 1687.430 1332.060 1687.750 ;
        RECT 1333.180 1687.430 1333.440 1687.750 ;
        RECT 1333.240 1684.010 1333.380 1687.430 ;
        RECT 1333.180 1683.690 1333.440 1684.010 ;
        RECT 1766.500 1674.170 1766.760 1674.490 ;
        RECT 1766.560 6.530 1766.700 1674.170 ;
        RECT 1766.560 6.390 1769.000 6.530 ;
        RECT 1768.860 2.400 1769.000 6.390 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1337.365 1661.325 1337.535 1687.675 ;
      LAYER mcon ;
        RECT 1337.365 1687.505 1337.535 1687.675 ;
      LAYER met1 ;
        RECT 1333.610 1687.660 1333.930 1687.720 ;
        RECT 1337.305 1687.660 1337.595 1687.705 ;
        RECT 1333.610 1687.520 1337.595 1687.660 ;
        RECT 1333.610 1687.460 1333.930 1687.520 ;
        RECT 1337.305 1687.475 1337.595 1687.520 ;
        RECT 1337.305 1661.480 1337.595 1661.525 ;
        RECT 1337.305 1661.340 1359.140 1661.480 ;
        RECT 1337.305 1661.295 1337.595 1661.340 ;
        RECT 1359.000 1660.800 1359.140 1661.340 ;
        RECT 1780.270 1660.800 1780.590 1660.860 ;
        RECT 1359.000 1660.660 1780.590 1660.800 ;
        RECT 1780.270 1660.600 1780.590 1660.660 ;
        RECT 1780.270 20.980 1780.590 21.040 ;
        RECT 1786.710 20.980 1787.030 21.040 ;
        RECT 1780.270 20.840 1787.030 20.980 ;
        RECT 1780.270 20.780 1780.590 20.840 ;
        RECT 1786.710 20.780 1787.030 20.840 ;
      LAYER via ;
        RECT 1333.640 1687.460 1333.900 1687.720 ;
        RECT 1780.300 1660.600 1780.560 1660.860 ;
        RECT 1780.300 20.780 1780.560 21.040 ;
        RECT 1786.740 20.780 1787.000 21.040 ;
      LAYER met2 ;
        RECT 1333.540 1700.340 1333.820 1704.000 ;
        RECT 1333.540 1700.000 1333.840 1700.340 ;
        RECT 1333.700 1687.750 1333.840 1700.000 ;
        RECT 1333.640 1687.430 1333.900 1687.750 ;
        RECT 1780.300 1660.570 1780.560 1660.890 ;
        RECT 1780.360 21.070 1780.500 1660.570 ;
        RECT 1780.300 20.750 1780.560 21.070 ;
        RECT 1786.740 20.750 1787.000 21.070 ;
        RECT 1786.800 2.400 1786.940 20.750 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1331.770 1676.780 1332.090 1676.840 ;
        RECT 1334.990 1676.780 1335.310 1676.840 ;
        RECT 1331.770 1676.640 1335.310 1676.780 ;
        RECT 1331.770 1676.580 1332.090 1676.640 ;
        RECT 1334.990 1676.580 1335.310 1676.640 ;
        RECT 1331.770 1633.260 1332.090 1633.320 ;
        RECT 1800.970 1633.260 1801.290 1633.320 ;
        RECT 1331.770 1633.120 1801.290 1633.260 ;
        RECT 1331.770 1633.060 1332.090 1633.120 ;
        RECT 1800.970 1633.060 1801.290 1633.120 ;
      LAYER via ;
        RECT 1331.800 1676.580 1332.060 1676.840 ;
        RECT 1335.020 1676.580 1335.280 1676.840 ;
        RECT 1331.800 1633.060 1332.060 1633.320 ;
        RECT 1801.000 1633.060 1801.260 1633.320 ;
      LAYER met2 ;
        RECT 1335.380 1700.410 1335.660 1704.000 ;
        RECT 1335.080 1700.270 1335.660 1700.410 ;
        RECT 1335.080 1676.870 1335.220 1700.270 ;
        RECT 1335.380 1700.000 1335.660 1700.270 ;
        RECT 1331.800 1676.550 1332.060 1676.870 ;
        RECT 1335.020 1676.550 1335.280 1676.870 ;
        RECT 1331.860 1633.350 1332.000 1676.550 ;
        RECT 1331.800 1633.030 1332.060 1633.350 ;
        RECT 1801.000 1633.030 1801.260 1633.350 ;
        RECT 1801.060 17.410 1801.200 1633.030 ;
        RECT 1801.060 17.270 1804.880 17.410 ;
        RECT 1804.740 2.400 1804.880 17.270 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1335.450 1684.260 1335.770 1684.320 ;
        RECT 1337.290 1684.260 1337.610 1684.320 ;
        RECT 1335.450 1684.120 1337.610 1684.260 ;
        RECT 1335.450 1684.060 1335.770 1684.120 ;
        RECT 1337.290 1684.060 1337.610 1684.120 ;
        RECT 1335.450 1598.240 1335.770 1598.300 ;
        RECT 1821.670 1598.240 1821.990 1598.300 ;
        RECT 1335.450 1598.100 1821.990 1598.240 ;
        RECT 1335.450 1598.040 1335.770 1598.100 ;
        RECT 1821.670 1598.040 1821.990 1598.100 ;
      LAYER via ;
        RECT 1335.480 1684.060 1335.740 1684.320 ;
        RECT 1337.320 1684.060 1337.580 1684.320 ;
        RECT 1335.480 1598.040 1335.740 1598.300 ;
        RECT 1821.700 1598.040 1821.960 1598.300 ;
      LAYER met2 ;
        RECT 1337.220 1700.340 1337.500 1704.000 ;
        RECT 1337.220 1700.000 1337.520 1700.340 ;
        RECT 1337.380 1684.350 1337.520 1700.000 ;
        RECT 1335.480 1684.030 1335.740 1684.350 ;
        RECT 1337.320 1684.030 1337.580 1684.350 ;
        RECT 1335.540 1598.330 1335.680 1684.030 ;
        RECT 1335.480 1598.010 1335.740 1598.330 ;
        RECT 1821.700 1598.010 1821.960 1598.330 ;
        RECT 1821.760 17.410 1821.900 1598.010 ;
        RECT 1821.760 17.270 1822.820 17.410 ;
        RECT 1822.680 2.400 1822.820 17.270 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1339.130 1684.260 1339.450 1684.320 ;
        RECT 1341.890 1684.260 1342.210 1684.320 ;
        RECT 1339.130 1684.120 1342.210 1684.260 ;
        RECT 1339.130 1684.060 1339.450 1684.120 ;
        RECT 1341.890 1684.060 1342.210 1684.120 ;
        RECT 1341.890 1626.120 1342.210 1626.180 ;
        RECT 1835.470 1626.120 1835.790 1626.180 ;
        RECT 1341.890 1625.980 1835.790 1626.120 ;
        RECT 1341.890 1625.920 1342.210 1625.980 ;
        RECT 1835.470 1625.920 1835.790 1625.980 ;
      LAYER via ;
        RECT 1339.160 1684.060 1339.420 1684.320 ;
        RECT 1341.920 1684.060 1342.180 1684.320 ;
        RECT 1341.920 1625.920 1342.180 1626.180 ;
        RECT 1835.500 1625.920 1835.760 1626.180 ;
      LAYER met2 ;
        RECT 1339.060 1700.340 1339.340 1704.000 ;
        RECT 1339.060 1700.000 1339.360 1700.340 ;
        RECT 1339.220 1684.350 1339.360 1700.000 ;
        RECT 1339.160 1684.030 1339.420 1684.350 ;
        RECT 1341.920 1684.030 1342.180 1684.350 ;
        RECT 1341.980 1626.210 1342.120 1684.030 ;
        RECT 1341.920 1625.890 1342.180 1626.210 ;
        RECT 1835.500 1625.890 1835.760 1626.210 ;
        RECT 1835.560 17.410 1835.700 1625.890 ;
        RECT 1835.560 17.270 1840.300 17.410 ;
        RECT 1840.160 2.400 1840.300 17.270 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1341.430 1584.640 1341.750 1584.700 ;
        RECT 1856.170 1584.640 1856.490 1584.700 ;
        RECT 1341.430 1584.500 1856.490 1584.640 ;
        RECT 1341.430 1584.440 1341.750 1584.500 ;
        RECT 1856.170 1584.440 1856.490 1584.500 ;
      LAYER via ;
        RECT 1341.460 1584.440 1341.720 1584.700 ;
        RECT 1856.200 1584.440 1856.460 1584.700 ;
      LAYER met2 ;
        RECT 1340.900 1700.340 1341.180 1704.000 ;
        RECT 1340.900 1700.000 1341.200 1700.340 ;
        RECT 1341.060 1661.140 1341.200 1700.000 ;
        RECT 1341.060 1661.000 1341.660 1661.140 ;
        RECT 1341.520 1584.730 1341.660 1661.000 ;
        RECT 1341.460 1584.410 1341.720 1584.730 ;
        RECT 1856.200 1584.410 1856.460 1584.730 ;
        RECT 1856.260 17.410 1856.400 1584.410 ;
        RECT 1856.260 17.270 1858.240 17.410 ;
        RECT 1858.100 2.400 1858.240 17.270 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1342.810 1678.480 1343.130 1678.540 ;
        RECT 1344.650 1678.480 1344.970 1678.540 ;
        RECT 1342.810 1678.340 1344.970 1678.480 ;
        RECT 1342.810 1678.280 1343.130 1678.340 ;
        RECT 1344.650 1678.280 1344.970 1678.340 ;
        RECT 1344.650 1667.600 1344.970 1667.660 ;
        RECT 1869.970 1667.600 1870.290 1667.660 ;
        RECT 1344.650 1667.460 1870.290 1667.600 ;
        RECT 1344.650 1667.400 1344.970 1667.460 ;
        RECT 1869.970 1667.400 1870.290 1667.460 ;
        RECT 1869.970 20.980 1870.290 21.040 ;
        RECT 1875.950 20.980 1876.270 21.040 ;
        RECT 1869.970 20.840 1876.270 20.980 ;
        RECT 1869.970 20.780 1870.290 20.840 ;
        RECT 1875.950 20.780 1876.270 20.840 ;
      LAYER via ;
        RECT 1342.840 1678.280 1343.100 1678.540 ;
        RECT 1344.680 1678.280 1344.940 1678.540 ;
        RECT 1344.680 1667.400 1344.940 1667.660 ;
        RECT 1870.000 1667.400 1870.260 1667.660 ;
        RECT 1870.000 20.780 1870.260 21.040 ;
        RECT 1875.980 20.780 1876.240 21.040 ;
      LAYER met2 ;
        RECT 1342.740 1700.340 1343.020 1704.000 ;
        RECT 1342.740 1700.000 1343.040 1700.340 ;
        RECT 1342.900 1678.570 1343.040 1700.000 ;
        RECT 1342.840 1678.250 1343.100 1678.570 ;
        RECT 1344.680 1678.250 1344.940 1678.570 ;
        RECT 1344.740 1667.690 1344.880 1678.250 ;
        RECT 1344.680 1667.370 1344.940 1667.690 ;
        RECT 1870.000 1667.370 1870.260 1667.690 ;
        RECT 1870.060 21.070 1870.200 1667.370 ;
        RECT 1870.000 20.750 1870.260 21.070 ;
        RECT 1875.980 20.750 1876.240 21.070 ;
        RECT 1876.040 2.400 1876.180 20.750 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1226.045 1601.485 1226.215 1642.115 ;
        RECT 1226.045 1558.985 1226.215 1593.835 ;
        RECT 1225.125 855.525 1225.295 903.975 ;
        RECT 1225.125 758.965 1225.295 807.075 ;
        RECT 1226.045 675.665 1226.215 693.515 ;
        RECT 1225.585 572.645 1225.755 620.755 ;
        RECT 1226.045 379.525 1226.215 427.635 ;
        RECT 1225.585 338.045 1225.755 352.495 ;
        RECT 1226.045 241.485 1226.215 289.595 ;
      LAYER mcon ;
        RECT 1226.045 1641.945 1226.215 1642.115 ;
        RECT 1226.045 1593.665 1226.215 1593.835 ;
        RECT 1225.125 903.805 1225.295 903.975 ;
        RECT 1225.125 806.905 1225.295 807.075 ;
        RECT 1226.045 693.345 1226.215 693.515 ;
        RECT 1225.585 620.585 1225.755 620.755 ;
        RECT 1226.045 427.465 1226.215 427.635 ;
        RECT 1225.585 352.325 1225.755 352.495 ;
        RECT 1226.045 289.425 1226.215 289.595 ;
      LAYER met1 ;
        RECT 1225.985 1642.100 1226.275 1642.145 ;
        RECT 1226.890 1642.100 1227.210 1642.160 ;
        RECT 1225.985 1641.960 1227.210 1642.100 ;
        RECT 1225.985 1641.915 1226.275 1641.960 ;
        RECT 1226.890 1641.900 1227.210 1641.960 ;
        RECT 1225.970 1601.640 1226.290 1601.700 ;
        RECT 1225.775 1601.500 1226.290 1601.640 ;
        RECT 1225.970 1601.440 1226.290 1601.500 ;
        RECT 1225.970 1593.820 1226.290 1593.880 ;
        RECT 1225.775 1593.680 1226.290 1593.820 ;
        RECT 1225.970 1593.620 1226.290 1593.680 ;
        RECT 1225.970 1559.140 1226.290 1559.200 ;
        RECT 1225.775 1559.000 1226.290 1559.140 ;
        RECT 1225.970 1558.940 1226.290 1559.000 ;
        RECT 1225.050 1062.740 1225.370 1062.800 ;
        RECT 1225.970 1062.740 1226.290 1062.800 ;
        RECT 1225.050 1062.600 1226.290 1062.740 ;
        RECT 1225.050 1062.540 1225.370 1062.600 ;
        RECT 1225.970 1062.540 1226.290 1062.600 ;
        RECT 1225.050 966.180 1225.370 966.240 ;
        RECT 1225.970 966.180 1226.290 966.240 ;
        RECT 1225.050 966.040 1226.290 966.180 ;
        RECT 1225.050 965.980 1225.370 966.040 ;
        RECT 1225.970 965.980 1226.290 966.040 ;
        RECT 1225.050 903.960 1225.370 904.020 ;
        RECT 1224.855 903.820 1225.370 903.960 ;
        RECT 1225.050 903.760 1225.370 903.820 ;
        RECT 1225.065 855.680 1225.355 855.725 ;
        RECT 1226.430 855.680 1226.750 855.740 ;
        RECT 1225.065 855.540 1226.750 855.680 ;
        RECT 1225.065 855.495 1225.355 855.540 ;
        RECT 1226.430 855.480 1226.750 855.540 ;
        RECT 1225.065 807.060 1225.355 807.105 ;
        RECT 1226.430 807.060 1226.750 807.120 ;
        RECT 1225.065 806.920 1226.750 807.060 ;
        RECT 1225.065 806.875 1225.355 806.920 ;
        RECT 1226.430 806.860 1226.750 806.920 ;
        RECT 1225.050 759.120 1225.370 759.180 ;
        RECT 1224.855 758.980 1225.370 759.120 ;
        RECT 1225.050 758.920 1225.370 758.980 ;
        RECT 1225.970 693.500 1226.290 693.560 ;
        RECT 1225.775 693.360 1226.290 693.500 ;
        RECT 1225.970 693.300 1226.290 693.360 ;
        RECT 1225.985 675.820 1226.275 675.865 ;
        RECT 1226.890 675.820 1227.210 675.880 ;
        RECT 1225.985 675.680 1227.210 675.820 ;
        RECT 1225.985 675.635 1226.275 675.680 ;
        RECT 1226.890 675.620 1227.210 675.680 ;
        RECT 1225.510 627.540 1225.830 627.600 ;
        RECT 1226.890 627.540 1227.210 627.600 ;
        RECT 1225.510 627.400 1227.210 627.540 ;
        RECT 1225.510 627.340 1225.830 627.400 ;
        RECT 1226.890 627.340 1227.210 627.400 ;
        RECT 1225.510 620.740 1225.830 620.800 ;
        RECT 1225.315 620.600 1225.830 620.740 ;
        RECT 1225.510 620.540 1225.830 620.600 ;
        RECT 1225.510 572.800 1225.830 572.860 ;
        RECT 1225.315 572.660 1225.830 572.800 ;
        RECT 1225.510 572.600 1225.830 572.660 ;
        RECT 1225.510 545.060 1225.830 545.320 ;
        RECT 1225.600 544.920 1225.740 545.060 ;
        RECT 1225.970 544.920 1226.290 544.980 ;
        RECT 1225.600 544.780 1226.290 544.920 ;
        RECT 1225.970 544.720 1226.290 544.780 ;
        RECT 1225.970 427.620 1226.290 427.680 ;
        RECT 1225.775 427.480 1226.290 427.620 ;
        RECT 1225.970 427.420 1226.290 427.480 ;
        RECT 1225.970 379.680 1226.290 379.740 ;
        RECT 1225.775 379.540 1226.290 379.680 ;
        RECT 1225.970 379.480 1226.290 379.540 ;
        RECT 1225.525 352.480 1225.815 352.525 ;
        RECT 1225.970 352.480 1226.290 352.540 ;
        RECT 1225.525 352.340 1226.290 352.480 ;
        RECT 1225.525 352.295 1225.815 352.340 ;
        RECT 1225.970 352.280 1226.290 352.340 ;
        RECT 1225.510 338.200 1225.830 338.260 ;
        RECT 1225.315 338.060 1225.830 338.200 ;
        RECT 1225.510 338.000 1225.830 338.060 ;
        RECT 1225.985 289.580 1226.275 289.625 ;
        RECT 1226.430 289.580 1226.750 289.640 ;
        RECT 1225.985 289.440 1226.750 289.580 ;
        RECT 1225.985 289.395 1226.275 289.440 ;
        RECT 1226.430 289.380 1226.750 289.440 ;
        RECT 1225.970 241.640 1226.290 241.700 ;
        RECT 1225.775 241.500 1226.290 241.640 ;
        RECT 1225.970 241.440 1226.290 241.500 ;
        RECT 758.150 79.460 758.470 79.520 ;
        RECT 1226.430 79.460 1226.750 79.520 ;
        RECT 758.150 79.320 1226.750 79.460 ;
        RECT 758.150 79.260 758.470 79.320 ;
        RECT 1226.430 79.260 1226.750 79.320 ;
        RECT 752.170 20.980 752.490 21.040 ;
        RECT 758.150 20.980 758.470 21.040 ;
        RECT 752.170 20.840 758.470 20.980 ;
        RECT 752.170 20.780 752.490 20.840 ;
        RECT 758.150 20.780 758.470 20.840 ;
      LAYER via ;
        RECT 1226.920 1641.900 1227.180 1642.160 ;
        RECT 1226.000 1601.440 1226.260 1601.700 ;
        RECT 1226.000 1593.620 1226.260 1593.880 ;
        RECT 1226.000 1558.940 1226.260 1559.200 ;
        RECT 1225.080 1062.540 1225.340 1062.800 ;
        RECT 1226.000 1062.540 1226.260 1062.800 ;
        RECT 1225.080 965.980 1225.340 966.240 ;
        RECT 1226.000 965.980 1226.260 966.240 ;
        RECT 1225.080 903.760 1225.340 904.020 ;
        RECT 1226.460 855.480 1226.720 855.740 ;
        RECT 1226.460 806.860 1226.720 807.120 ;
        RECT 1225.080 758.920 1225.340 759.180 ;
        RECT 1226.000 693.300 1226.260 693.560 ;
        RECT 1226.920 675.620 1227.180 675.880 ;
        RECT 1225.540 627.340 1225.800 627.600 ;
        RECT 1226.920 627.340 1227.180 627.600 ;
        RECT 1225.540 620.540 1225.800 620.800 ;
        RECT 1225.540 572.600 1225.800 572.860 ;
        RECT 1225.540 545.060 1225.800 545.320 ;
        RECT 1226.000 544.720 1226.260 544.980 ;
        RECT 1226.000 427.420 1226.260 427.680 ;
        RECT 1226.000 379.480 1226.260 379.740 ;
        RECT 1226.000 352.280 1226.260 352.540 ;
        RECT 1225.540 338.000 1225.800 338.260 ;
        RECT 1226.460 289.380 1226.720 289.640 ;
        RECT 1226.000 241.440 1226.260 241.700 ;
        RECT 758.180 79.260 758.440 79.520 ;
        RECT 1226.460 79.260 1226.720 79.520 ;
        RECT 752.200 20.780 752.460 21.040 ;
        RECT 758.180 20.780 758.440 21.040 ;
      LAYER met2 ;
        RECT 1226.820 1700.340 1227.100 1704.000 ;
        RECT 1226.820 1700.000 1227.120 1700.340 ;
        RECT 1226.980 1642.190 1227.120 1700.000 ;
        RECT 1226.920 1641.870 1227.180 1642.190 ;
        RECT 1226.000 1601.410 1226.260 1601.730 ;
        RECT 1226.060 1593.910 1226.200 1601.410 ;
        RECT 1226.000 1593.590 1226.260 1593.910 ;
        RECT 1226.000 1558.910 1226.260 1559.230 ;
        RECT 1226.060 1125.130 1226.200 1558.910 ;
        RECT 1225.600 1124.990 1226.200 1125.130 ;
        RECT 1225.600 1124.450 1225.740 1124.990 ;
        RECT 1225.600 1124.310 1226.200 1124.450 ;
        RECT 1226.060 1110.965 1226.200 1124.310 ;
        RECT 1225.070 1110.595 1225.350 1110.965 ;
        RECT 1225.990 1110.595 1226.270 1110.965 ;
        RECT 1225.140 1062.830 1225.280 1110.595 ;
        RECT 1225.080 1062.510 1225.340 1062.830 ;
        RECT 1226.000 1062.510 1226.260 1062.830 ;
        RECT 1226.060 1014.405 1226.200 1062.510 ;
        RECT 1225.070 1014.035 1225.350 1014.405 ;
        RECT 1225.990 1014.035 1226.270 1014.405 ;
        RECT 1225.140 966.270 1225.280 1014.035 ;
        RECT 1225.080 965.950 1225.340 966.270 ;
        RECT 1226.000 965.950 1226.260 966.270 ;
        RECT 1226.060 917.845 1226.200 965.950 ;
        RECT 1225.070 917.475 1225.350 917.845 ;
        RECT 1225.990 917.475 1226.270 917.845 ;
        RECT 1225.140 904.050 1225.280 917.475 ;
        RECT 1225.080 903.730 1225.340 904.050 ;
        RECT 1226.460 855.450 1226.720 855.770 ;
        RECT 1226.520 807.150 1226.660 855.450 ;
        RECT 1226.460 806.830 1226.720 807.150 ;
        RECT 1225.080 758.890 1225.340 759.210 ;
        RECT 1225.140 717.925 1225.280 758.890 ;
        RECT 1225.070 717.555 1225.350 717.925 ;
        RECT 1225.990 717.555 1226.270 717.925 ;
        RECT 1226.060 693.590 1226.200 717.555 ;
        RECT 1226.000 693.270 1226.260 693.590 ;
        RECT 1226.920 675.590 1227.180 675.910 ;
        RECT 1226.980 669.530 1227.120 675.590 ;
        RECT 1226.980 669.390 1227.580 669.530 ;
        RECT 1227.440 641.650 1227.580 669.390 ;
        RECT 1226.980 641.510 1227.580 641.650 ;
        RECT 1226.980 627.630 1227.120 641.510 ;
        RECT 1225.540 627.310 1225.800 627.630 ;
        RECT 1226.920 627.310 1227.180 627.630 ;
        RECT 1225.600 620.830 1225.740 627.310 ;
        RECT 1225.540 620.510 1225.800 620.830 ;
        RECT 1225.540 572.570 1225.800 572.890 ;
        RECT 1225.600 545.350 1225.740 572.570 ;
        RECT 1225.540 545.030 1225.800 545.350 ;
        RECT 1226.000 544.690 1226.260 545.010 ;
        RECT 1226.060 530.810 1226.200 544.690 ;
        RECT 1226.060 530.670 1226.660 530.810 ;
        RECT 1226.520 448.530 1226.660 530.670 ;
        RECT 1226.060 448.390 1226.660 448.530 ;
        RECT 1226.060 427.710 1226.200 448.390 ;
        RECT 1226.000 427.390 1226.260 427.710 ;
        RECT 1226.000 379.450 1226.260 379.770 ;
        RECT 1226.060 352.570 1226.200 379.450 ;
        RECT 1226.000 352.250 1226.260 352.570 ;
        RECT 1225.540 337.970 1225.800 338.290 ;
        RECT 1225.600 324.770 1225.740 337.970 ;
        RECT 1225.600 324.630 1226.660 324.770 ;
        RECT 1226.520 289.670 1226.660 324.630 ;
        RECT 1226.460 289.350 1226.720 289.670 ;
        RECT 1226.000 241.410 1226.260 241.730 ;
        RECT 1226.060 207.130 1226.200 241.410 ;
        RECT 1226.060 206.990 1226.660 207.130 ;
        RECT 1226.520 79.550 1226.660 206.990 ;
        RECT 758.180 79.230 758.440 79.550 ;
        RECT 1226.460 79.230 1226.720 79.550 ;
        RECT 758.240 21.070 758.380 79.230 ;
        RECT 752.200 20.750 752.460 21.070 ;
        RECT 758.180 20.750 758.440 21.070 ;
        RECT 752.260 2.400 752.400 20.750 ;
        RECT 752.050 -4.800 752.610 2.400 ;
      LAYER via2 ;
        RECT 1225.070 1110.640 1225.350 1110.920 ;
        RECT 1225.990 1110.640 1226.270 1110.920 ;
        RECT 1225.070 1014.080 1225.350 1014.360 ;
        RECT 1225.990 1014.080 1226.270 1014.360 ;
        RECT 1225.070 917.520 1225.350 917.800 ;
        RECT 1225.990 917.520 1226.270 917.800 ;
        RECT 1225.070 717.600 1225.350 717.880 ;
        RECT 1225.990 717.600 1226.270 717.880 ;
      LAYER met3 ;
        RECT 1225.045 1110.930 1225.375 1110.945 ;
        RECT 1225.965 1110.930 1226.295 1110.945 ;
        RECT 1225.045 1110.630 1226.295 1110.930 ;
        RECT 1225.045 1110.615 1225.375 1110.630 ;
        RECT 1225.965 1110.615 1226.295 1110.630 ;
        RECT 1225.045 1014.370 1225.375 1014.385 ;
        RECT 1225.965 1014.370 1226.295 1014.385 ;
        RECT 1225.045 1014.070 1226.295 1014.370 ;
        RECT 1225.045 1014.055 1225.375 1014.070 ;
        RECT 1225.965 1014.055 1226.295 1014.070 ;
        RECT 1225.045 917.810 1225.375 917.825 ;
        RECT 1225.965 917.810 1226.295 917.825 ;
        RECT 1225.045 917.510 1226.295 917.810 ;
        RECT 1225.045 917.495 1225.375 917.510 ;
        RECT 1225.965 917.495 1226.295 917.510 ;
        RECT 1225.045 717.890 1225.375 717.905 ;
        RECT 1225.965 717.890 1226.295 717.905 ;
        RECT 1225.045 717.590 1226.295 717.890 ;
        RECT 1225.045 717.575 1225.375 717.590 ;
        RECT 1225.965 717.575 1226.295 717.590 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1342.810 1677.460 1343.130 1677.520 ;
        RECT 1344.190 1677.460 1344.510 1677.520 ;
        RECT 1342.810 1677.320 1344.510 1677.460 ;
        RECT 1342.810 1677.260 1343.130 1677.320 ;
        RECT 1344.190 1677.260 1344.510 1677.320 ;
        RECT 1342.810 1556.420 1343.130 1556.480 ;
        RECT 1890.670 1556.420 1890.990 1556.480 ;
        RECT 1342.810 1556.280 1890.990 1556.420 ;
        RECT 1342.810 1556.220 1343.130 1556.280 ;
        RECT 1890.670 1556.220 1890.990 1556.280 ;
      LAYER via ;
        RECT 1342.840 1677.260 1343.100 1677.520 ;
        RECT 1344.220 1677.260 1344.480 1677.520 ;
        RECT 1342.840 1556.220 1343.100 1556.480 ;
        RECT 1890.700 1556.220 1890.960 1556.480 ;
      LAYER met2 ;
        RECT 1344.580 1700.410 1344.860 1704.000 ;
        RECT 1344.280 1700.270 1344.860 1700.410 ;
        RECT 1344.280 1677.550 1344.420 1700.270 ;
        RECT 1344.580 1700.000 1344.860 1700.270 ;
        RECT 1342.840 1677.230 1343.100 1677.550 ;
        RECT 1344.220 1677.230 1344.480 1677.550 ;
        RECT 1342.900 1556.510 1343.040 1677.230 ;
        RECT 1342.840 1556.190 1343.100 1556.510 ;
        RECT 1890.700 1556.190 1890.960 1556.510 ;
        RECT 1890.760 17.410 1890.900 1556.190 ;
        RECT 1890.760 17.270 1894.120 17.410 ;
        RECT 1893.980 2.400 1894.120 17.270 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.490 1640.060 1346.810 1640.120 ;
        RECT 1911.370 1640.060 1911.690 1640.120 ;
        RECT 1346.490 1639.920 1911.690 1640.060 ;
        RECT 1346.490 1639.860 1346.810 1639.920 ;
        RECT 1911.370 1639.860 1911.690 1639.920 ;
      LAYER via ;
        RECT 1346.520 1639.860 1346.780 1640.120 ;
        RECT 1911.400 1639.860 1911.660 1640.120 ;
      LAYER met2 ;
        RECT 1346.420 1700.340 1346.700 1704.000 ;
        RECT 1346.420 1700.000 1346.720 1700.340 ;
        RECT 1346.580 1640.150 1346.720 1700.000 ;
        RECT 1346.520 1639.830 1346.780 1640.150 ;
        RECT 1911.400 1639.830 1911.660 1640.150 ;
        RECT 1911.460 17.410 1911.600 1639.830 ;
        RECT 1911.460 17.270 1912.060 17.410 ;
        RECT 1911.920 2.400 1912.060 17.270 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1348.790 1619.320 1349.110 1619.380 ;
        RECT 1925.170 1619.320 1925.490 1619.380 ;
        RECT 1348.790 1619.180 1925.490 1619.320 ;
        RECT 1348.790 1619.120 1349.110 1619.180 ;
        RECT 1925.170 1619.120 1925.490 1619.180 ;
      LAYER via ;
        RECT 1348.820 1619.120 1349.080 1619.380 ;
        RECT 1925.200 1619.120 1925.460 1619.380 ;
      LAYER met2 ;
        RECT 1348.260 1700.340 1348.540 1704.000 ;
        RECT 1348.260 1700.000 1348.560 1700.340 ;
        RECT 1348.420 1635.130 1348.560 1700.000 ;
        RECT 1348.420 1634.990 1349.020 1635.130 ;
        RECT 1348.880 1619.410 1349.020 1634.990 ;
        RECT 1348.820 1619.090 1349.080 1619.410 ;
        RECT 1925.200 1619.090 1925.460 1619.410 ;
        RECT 1925.260 17.410 1925.400 1619.090 ;
        RECT 1925.260 17.270 1929.540 17.410 ;
        RECT 1929.400 2.400 1929.540 17.270 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1349.710 1549.620 1350.030 1549.680 ;
        RECT 1945.870 1549.620 1946.190 1549.680 ;
        RECT 1349.710 1549.480 1946.190 1549.620 ;
        RECT 1349.710 1549.420 1350.030 1549.480 ;
        RECT 1945.870 1549.420 1946.190 1549.480 ;
      LAYER via ;
        RECT 1349.740 1549.420 1350.000 1549.680 ;
        RECT 1945.900 1549.420 1946.160 1549.680 ;
      LAYER met2 ;
        RECT 1350.100 1700.410 1350.380 1704.000 ;
        RECT 1349.800 1700.270 1350.380 1700.410 ;
        RECT 1349.800 1549.710 1349.940 1700.270 ;
        RECT 1350.100 1700.000 1350.380 1700.270 ;
        RECT 1349.740 1549.390 1350.000 1549.710 ;
        RECT 1945.900 1549.390 1946.160 1549.710 ;
        RECT 1945.960 17.410 1946.100 1549.390 ;
        RECT 1945.960 17.270 1947.480 17.410 ;
        RECT 1947.340 2.400 1947.480 17.270 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1347.945 268.005 1348.115 282.795 ;
      LAYER mcon ;
        RECT 1347.945 282.625 1348.115 282.795 ;
      LAYER met1 ;
        RECT 1347.410 1678.140 1347.730 1678.200 ;
        RECT 1351.550 1678.140 1351.870 1678.200 ;
        RECT 1347.410 1678.000 1351.870 1678.140 ;
        RECT 1347.410 1677.940 1347.730 1678.000 ;
        RECT 1351.550 1677.940 1351.870 1678.000 ;
        RECT 1348.330 1539.420 1348.650 1539.480 ;
        RECT 1347.960 1539.280 1348.650 1539.420 ;
        RECT 1347.960 1538.460 1348.100 1539.280 ;
        RECT 1348.330 1539.220 1348.650 1539.280 ;
        RECT 1347.870 1538.200 1348.190 1538.460 ;
        RECT 1347.870 282.780 1348.190 282.840 ;
        RECT 1347.675 282.640 1348.190 282.780 ;
        RECT 1347.870 282.580 1348.190 282.640 ;
        RECT 1347.885 268.160 1348.175 268.205 ;
        RECT 1348.330 268.160 1348.650 268.220 ;
        RECT 1347.885 268.020 1348.650 268.160 ;
        RECT 1347.885 267.975 1348.175 268.020 ;
        RECT 1348.330 267.960 1348.650 268.020 ;
        RECT 1347.870 186.220 1348.190 186.280 ;
        RECT 1348.330 186.220 1348.650 186.280 ;
        RECT 1347.870 186.080 1348.650 186.220 ;
        RECT 1347.870 186.020 1348.190 186.080 ;
        RECT 1348.330 186.020 1348.650 186.080 ;
        RECT 1348.330 90.340 1348.650 90.400 ;
        RECT 1347.960 90.200 1348.650 90.340 ;
        RECT 1347.960 90.060 1348.100 90.200 ;
        RECT 1348.330 90.140 1348.650 90.200 ;
        RECT 1347.870 89.800 1348.190 90.060 ;
        RECT 1348.330 42.060 1348.650 42.120 ;
        RECT 1347.960 41.920 1348.650 42.060 ;
        RECT 1347.960 41.780 1348.100 41.920 ;
        RECT 1348.330 41.860 1348.650 41.920 ;
        RECT 1347.870 41.520 1348.190 41.780 ;
        RECT 1347.870 14.180 1348.190 14.240 ;
        RECT 1965.190 14.180 1965.510 14.240 ;
        RECT 1347.870 14.040 1952.540 14.180 ;
        RECT 1347.870 13.980 1348.190 14.040 ;
        RECT 1952.400 13.840 1952.540 14.040 ;
        RECT 1959.760 14.040 1965.510 14.180 ;
        RECT 1959.760 13.840 1959.900 14.040 ;
        RECT 1965.190 13.980 1965.510 14.040 ;
        RECT 1952.400 13.700 1959.900 13.840 ;
      LAYER via ;
        RECT 1347.440 1677.940 1347.700 1678.200 ;
        RECT 1351.580 1677.940 1351.840 1678.200 ;
        RECT 1348.360 1539.220 1348.620 1539.480 ;
        RECT 1347.900 1538.200 1348.160 1538.460 ;
        RECT 1347.900 282.580 1348.160 282.840 ;
        RECT 1348.360 267.960 1348.620 268.220 ;
        RECT 1347.900 186.020 1348.160 186.280 ;
        RECT 1348.360 186.020 1348.620 186.280 ;
        RECT 1348.360 90.140 1348.620 90.400 ;
        RECT 1347.900 89.800 1348.160 90.060 ;
        RECT 1348.360 41.860 1348.620 42.120 ;
        RECT 1347.900 41.520 1348.160 41.780 ;
        RECT 1347.900 13.980 1348.160 14.240 ;
        RECT 1965.220 13.980 1965.480 14.240 ;
      LAYER met2 ;
        RECT 1351.940 1700.410 1352.220 1704.000 ;
        RECT 1351.640 1700.270 1352.220 1700.410 ;
        RECT 1351.640 1678.230 1351.780 1700.270 ;
        RECT 1351.940 1700.000 1352.220 1700.270 ;
        RECT 1347.440 1677.910 1347.700 1678.230 ;
        RECT 1351.580 1677.910 1351.840 1678.230 ;
        RECT 1347.500 1634.450 1347.640 1677.910 ;
        RECT 1347.500 1634.310 1348.560 1634.450 ;
        RECT 1348.420 1539.510 1348.560 1634.310 ;
        RECT 1348.360 1539.190 1348.620 1539.510 ;
        RECT 1347.900 1538.170 1348.160 1538.490 ;
        RECT 1347.960 282.870 1348.100 1538.170 ;
        RECT 1347.900 282.550 1348.160 282.870 ;
        RECT 1348.360 267.930 1348.620 268.250 ;
        RECT 1348.420 186.310 1348.560 267.930 ;
        RECT 1347.900 185.990 1348.160 186.310 ;
        RECT 1348.360 185.990 1348.620 186.310 ;
        RECT 1347.960 137.770 1348.100 185.990 ;
        RECT 1347.960 137.630 1348.560 137.770 ;
        RECT 1348.420 90.430 1348.560 137.630 ;
        RECT 1348.360 90.110 1348.620 90.430 ;
        RECT 1347.900 89.770 1348.160 90.090 ;
        RECT 1347.960 89.490 1348.100 89.770 ;
        RECT 1347.960 89.350 1348.560 89.490 ;
        RECT 1348.420 42.150 1348.560 89.350 ;
        RECT 1348.360 41.830 1348.620 42.150 ;
        RECT 1347.900 41.490 1348.160 41.810 ;
        RECT 1347.960 14.270 1348.100 41.490 ;
        RECT 1347.900 13.950 1348.160 14.270 ;
        RECT 1965.220 13.950 1965.480 14.270 ;
        RECT 1965.280 2.400 1965.420 13.950 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1358.065 931.685 1358.235 979.795 ;
        RECT 1358.065 745.705 1358.235 800.275 ;
        RECT 1358.065 697.425 1358.235 745.195 ;
        RECT 1357.605 648.805 1357.775 696.915 ;
        RECT 1358.065 89.845 1358.235 186.235 ;
      LAYER mcon ;
        RECT 1358.065 979.625 1358.235 979.795 ;
        RECT 1358.065 800.105 1358.235 800.275 ;
        RECT 1358.065 745.025 1358.235 745.195 ;
        RECT 1357.605 696.745 1357.775 696.915 ;
        RECT 1358.065 186.065 1358.235 186.235 ;
      LAYER met1 ;
        RECT 1353.850 1670.660 1354.170 1670.720 ;
        RECT 1358.910 1670.660 1359.230 1670.720 ;
        RECT 1353.850 1670.520 1359.230 1670.660 ;
        RECT 1353.850 1670.460 1354.170 1670.520 ;
        RECT 1358.910 1670.460 1359.230 1670.520 ;
        RECT 1357.530 1228.320 1357.850 1228.380 ;
        RECT 1358.910 1228.320 1359.230 1228.380 ;
        RECT 1357.530 1228.180 1359.230 1228.320 ;
        RECT 1357.530 1228.120 1357.850 1228.180 ;
        RECT 1358.910 1228.120 1359.230 1228.180 ;
        RECT 1357.990 1187.180 1358.310 1187.240 ;
        RECT 1358.910 1187.180 1359.230 1187.240 ;
        RECT 1357.990 1187.040 1359.230 1187.180 ;
        RECT 1357.990 1186.980 1358.310 1187.040 ;
        RECT 1358.910 1186.980 1359.230 1187.040 ;
        RECT 1357.990 979.780 1358.310 979.840 ;
        RECT 1357.795 979.640 1358.310 979.780 ;
        RECT 1357.990 979.580 1358.310 979.640 ;
        RECT 1358.005 931.840 1358.295 931.885 ;
        RECT 1358.450 931.840 1358.770 931.900 ;
        RECT 1358.005 931.700 1358.770 931.840 ;
        RECT 1358.005 931.655 1358.295 931.700 ;
        RECT 1358.450 931.640 1358.770 931.700 ;
        RECT 1357.990 890.360 1358.310 890.420 ;
        RECT 1358.450 890.360 1358.770 890.420 ;
        RECT 1357.990 890.220 1358.770 890.360 ;
        RECT 1357.990 890.160 1358.310 890.220 ;
        RECT 1358.450 890.160 1358.770 890.220 ;
        RECT 1357.990 800.260 1358.310 800.320 ;
        RECT 1357.795 800.120 1358.310 800.260 ;
        RECT 1357.990 800.060 1358.310 800.120 ;
        RECT 1358.005 745.860 1358.295 745.905 ;
        RECT 1358.450 745.860 1358.770 745.920 ;
        RECT 1358.005 745.720 1358.770 745.860 ;
        RECT 1358.005 745.675 1358.295 745.720 ;
        RECT 1358.450 745.660 1358.770 745.720 ;
        RECT 1357.990 745.180 1358.310 745.240 ;
        RECT 1357.795 745.040 1358.310 745.180 ;
        RECT 1357.990 744.980 1358.310 745.040 ;
        RECT 1357.990 697.580 1358.310 697.640 ;
        RECT 1357.795 697.440 1358.310 697.580 ;
        RECT 1357.990 697.380 1358.310 697.440 ;
        RECT 1357.545 696.900 1357.835 696.945 ;
        RECT 1357.990 696.900 1358.310 696.960 ;
        RECT 1357.545 696.760 1358.310 696.900 ;
        RECT 1357.545 696.715 1357.835 696.760 ;
        RECT 1357.990 696.700 1358.310 696.760 ;
        RECT 1357.530 648.960 1357.850 649.020 ;
        RECT 1357.530 648.820 1358.045 648.960 ;
        RECT 1357.530 648.760 1357.850 648.820 ;
        RECT 1357.990 186.220 1358.310 186.280 ;
        RECT 1357.795 186.080 1358.310 186.220 ;
        RECT 1357.990 186.020 1358.310 186.080 ;
        RECT 1357.990 90.000 1358.310 90.060 ;
        RECT 1357.795 89.860 1358.310 90.000 ;
        RECT 1357.990 89.800 1358.310 89.860 ;
        RECT 1357.990 14.520 1358.310 14.580 ;
        RECT 1983.130 14.520 1983.450 14.580 ;
        RECT 1357.990 14.380 1983.450 14.520 ;
        RECT 1357.990 14.320 1358.310 14.380 ;
        RECT 1983.130 14.320 1983.450 14.380 ;
      LAYER via ;
        RECT 1353.880 1670.460 1354.140 1670.720 ;
        RECT 1358.940 1670.460 1359.200 1670.720 ;
        RECT 1357.560 1228.120 1357.820 1228.380 ;
        RECT 1358.940 1228.120 1359.200 1228.380 ;
        RECT 1358.020 1186.980 1358.280 1187.240 ;
        RECT 1358.940 1186.980 1359.200 1187.240 ;
        RECT 1358.020 979.580 1358.280 979.840 ;
        RECT 1358.480 931.640 1358.740 931.900 ;
        RECT 1358.020 890.160 1358.280 890.420 ;
        RECT 1358.480 890.160 1358.740 890.420 ;
        RECT 1358.020 800.060 1358.280 800.320 ;
        RECT 1358.480 745.660 1358.740 745.920 ;
        RECT 1358.020 744.980 1358.280 745.240 ;
        RECT 1358.020 697.380 1358.280 697.640 ;
        RECT 1358.020 696.700 1358.280 696.960 ;
        RECT 1357.560 648.760 1357.820 649.020 ;
        RECT 1358.020 186.020 1358.280 186.280 ;
        RECT 1358.020 89.800 1358.280 90.060 ;
        RECT 1358.020 14.320 1358.280 14.580 ;
        RECT 1983.160 14.320 1983.420 14.580 ;
      LAYER met2 ;
        RECT 1353.780 1700.340 1354.060 1704.000 ;
        RECT 1353.780 1700.000 1354.080 1700.340 ;
        RECT 1353.940 1670.750 1354.080 1700.000 ;
        RECT 1353.880 1670.430 1354.140 1670.750 ;
        RECT 1358.940 1670.430 1359.200 1670.750 ;
        RECT 1359.000 1476.805 1359.140 1670.430 ;
        RECT 1358.010 1476.435 1358.290 1476.805 ;
        RECT 1358.930 1476.435 1359.210 1476.805 ;
        RECT 1358.080 1252.290 1358.220 1476.435 ;
        RECT 1357.620 1252.150 1358.220 1252.290 ;
        RECT 1357.620 1228.410 1357.760 1252.150 ;
        RECT 1357.560 1228.090 1357.820 1228.410 ;
        RECT 1358.940 1228.090 1359.200 1228.410 ;
        RECT 1359.000 1187.270 1359.140 1228.090 ;
        RECT 1358.020 1186.950 1358.280 1187.270 ;
        RECT 1358.940 1186.950 1359.200 1187.270 ;
        RECT 1358.080 979.870 1358.220 1186.950 ;
        RECT 1358.020 979.550 1358.280 979.870 ;
        RECT 1358.480 931.610 1358.740 931.930 ;
        RECT 1358.540 890.450 1358.680 931.610 ;
        RECT 1358.020 890.130 1358.280 890.450 ;
        RECT 1358.480 890.130 1358.740 890.450 ;
        RECT 1358.080 800.350 1358.220 890.130 ;
        RECT 1358.020 800.030 1358.280 800.350 ;
        RECT 1358.480 745.690 1358.740 745.950 ;
        RECT 1358.080 745.630 1358.740 745.690 ;
        RECT 1358.080 745.550 1358.680 745.630 ;
        RECT 1358.080 745.270 1358.220 745.550 ;
        RECT 1358.020 744.950 1358.280 745.270 ;
        RECT 1358.020 697.350 1358.280 697.670 ;
        RECT 1358.080 696.990 1358.220 697.350 ;
        RECT 1358.020 696.670 1358.280 696.990 ;
        RECT 1357.560 648.730 1357.820 649.050 ;
        RECT 1357.620 631.450 1357.760 648.730 ;
        RECT 1357.620 631.310 1358.220 631.450 ;
        RECT 1358.080 186.310 1358.220 631.310 ;
        RECT 1358.020 185.990 1358.280 186.310 ;
        RECT 1358.020 89.770 1358.280 90.090 ;
        RECT 1358.080 14.610 1358.220 89.770 ;
        RECT 1358.020 14.290 1358.280 14.610 ;
        RECT 1983.160 14.290 1983.420 14.610 ;
        RECT 1983.220 2.400 1983.360 14.290 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
      LAYER via2 ;
        RECT 1358.010 1476.480 1358.290 1476.760 ;
        RECT 1358.930 1476.480 1359.210 1476.760 ;
      LAYER met3 ;
        RECT 1357.985 1476.770 1358.315 1476.785 ;
        RECT 1358.905 1476.770 1359.235 1476.785 ;
        RECT 1357.985 1476.470 1359.235 1476.770 ;
        RECT 1357.985 1476.455 1358.315 1476.470 ;
        RECT 1358.905 1476.455 1359.235 1476.470 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1355.230 14.860 1355.550 14.920 ;
        RECT 2001.070 14.860 2001.390 14.920 ;
        RECT 1355.230 14.720 2001.390 14.860 ;
        RECT 1355.230 14.660 1355.550 14.720 ;
        RECT 2001.070 14.660 2001.390 14.720 ;
      LAYER via ;
        RECT 1355.260 14.660 1355.520 14.920 ;
        RECT 2001.100 14.660 2001.360 14.920 ;
      LAYER met2 ;
        RECT 1355.620 1700.410 1355.900 1704.000 ;
        RECT 1355.320 1700.270 1355.900 1700.410 ;
        RECT 1355.320 14.950 1355.460 1700.270 ;
        RECT 1355.620 1700.000 1355.900 1700.270 ;
        RECT 1355.260 14.630 1355.520 14.950 ;
        RECT 2001.100 14.630 2001.360 14.950 ;
        RECT 2001.160 2.400 2001.300 14.630 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1355.690 1497.600 1356.010 1497.660 ;
        RECT 1357.530 1497.600 1357.850 1497.660 ;
        RECT 1355.690 1497.460 1357.850 1497.600 ;
        RECT 1355.690 1497.400 1356.010 1497.460 ;
        RECT 1357.530 1497.400 1357.850 1497.460 ;
        RECT 1355.690 331.060 1356.010 331.120 ;
        RECT 1356.150 331.060 1356.470 331.120 ;
        RECT 1355.690 330.920 1356.470 331.060 ;
        RECT 1355.690 330.860 1356.010 330.920 ;
        RECT 1356.150 330.860 1356.470 330.920 ;
        RECT 1355.690 241.640 1356.010 241.700 ;
        RECT 1356.150 241.640 1356.470 241.700 ;
        RECT 1355.690 241.500 1356.470 241.640 ;
        RECT 1355.690 241.440 1356.010 241.500 ;
        RECT 1356.150 241.440 1356.470 241.500 ;
        RECT 1355.690 15.200 1356.010 15.260 ;
        RECT 2018.550 15.200 2018.870 15.260 ;
        RECT 1355.690 15.060 2018.870 15.200 ;
        RECT 1355.690 15.000 1356.010 15.060 ;
        RECT 2018.550 15.000 2018.870 15.060 ;
      LAYER via ;
        RECT 1355.720 1497.400 1355.980 1497.660 ;
        RECT 1357.560 1497.400 1357.820 1497.660 ;
        RECT 1355.720 330.860 1355.980 331.120 ;
        RECT 1356.180 330.860 1356.440 331.120 ;
        RECT 1355.720 241.440 1355.980 241.700 ;
        RECT 1356.180 241.440 1356.440 241.700 ;
        RECT 1355.720 15.000 1355.980 15.260 ;
        RECT 2018.580 15.000 2018.840 15.260 ;
      LAYER met2 ;
        RECT 1357.460 1700.340 1357.740 1704.000 ;
        RECT 1357.460 1700.000 1357.760 1700.340 ;
        RECT 1357.620 1497.690 1357.760 1700.000 ;
        RECT 1355.720 1497.370 1355.980 1497.690 ;
        RECT 1357.560 1497.370 1357.820 1497.690 ;
        RECT 1355.780 331.150 1355.920 1497.370 ;
        RECT 1355.720 330.830 1355.980 331.150 ;
        RECT 1356.180 330.830 1356.440 331.150 ;
        RECT 1356.240 241.730 1356.380 330.830 ;
        RECT 1355.720 241.410 1355.980 241.730 ;
        RECT 1356.180 241.410 1356.440 241.730 ;
        RECT 1355.780 15.290 1355.920 241.410 ;
        RECT 1355.720 14.970 1355.980 15.290 ;
        RECT 2018.580 14.970 2018.840 15.290 ;
        RECT 2018.640 2.400 2018.780 14.970 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1359.370 1666.580 1359.690 1666.640 ;
        RECT 1361.210 1666.580 1361.530 1666.640 ;
        RECT 1359.370 1666.440 1361.530 1666.580 ;
        RECT 1359.370 1666.380 1359.690 1666.440 ;
        RECT 1361.210 1666.380 1361.530 1666.440 ;
        RECT 1361.210 15.540 1361.530 15.600 ;
        RECT 2036.490 15.540 2036.810 15.600 ;
        RECT 1361.210 15.400 2036.810 15.540 ;
        RECT 1361.210 15.340 1361.530 15.400 ;
        RECT 2036.490 15.340 2036.810 15.400 ;
      LAYER via ;
        RECT 1359.400 1666.380 1359.660 1666.640 ;
        RECT 1361.240 1666.380 1361.500 1666.640 ;
        RECT 1361.240 15.340 1361.500 15.600 ;
        RECT 2036.520 15.340 2036.780 15.600 ;
      LAYER met2 ;
        RECT 1359.300 1700.340 1359.580 1704.000 ;
        RECT 1359.300 1700.000 1359.600 1700.340 ;
        RECT 1359.460 1666.670 1359.600 1700.000 ;
        RECT 1359.400 1666.350 1359.660 1666.670 ;
        RECT 1361.240 1666.350 1361.500 1666.670 ;
        RECT 1361.300 15.630 1361.440 1666.350 ;
        RECT 1361.240 15.310 1361.500 15.630 ;
        RECT 2036.520 15.310 2036.780 15.630 ;
        RECT 2036.580 2.400 2036.720 15.310 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1359.830 1683.920 1360.150 1683.980 ;
        RECT 1361.210 1683.920 1361.530 1683.980 ;
        RECT 1359.830 1683.780 1361.530 1683.920 ;
        RECT 1359.830 1683.720 1360.150 1683.780 ;
        RECT 1361.210 1683.720 1361.530 1683.780 ;
        RECT 1359.830 15.880 1360.150 15.940 ;
        RECT 2054.430 15.880 2054.750 15.940 ;
        RECT 1359.830 15.740 2054.750 15.880 ;
        RECT 1359.830 15.680 1360.150 15.740 ;
        RECT 2054.430 15.680 2054.750 15.740 ;
      LAYER via ;
        RECT 1359.860 1683.720 1360.120 1683.980 ;
        RECT 1361.240 1683.720 1361.500 1683.980 ;
        RECT 1359.860 15.680 1360.120 15.940 ;
        RECT 2054.460 15.680 2054.720 15.940 ;
      LAYER met2 ;
        RECT 1361.140 1700.340 1361.420 1704.000 ;
        RECT 1361.140 1700.000 1361.440 1700.340 ;
        RECT 1361.300 1684.010 1361.440 1700.000 ;
        RECT 1359.860 1683.690 1360.120 1684.010 ;
        RECT 1361.240 1683.690 1361.500 1684.010 ;
        RECT 1359.920 15.970 1360.060 1683.690 ;
        RECT 1359.860 15.650 1360.120 15.970 ;
        RECT 2054.460 15.650 2054.720 15.970 ;
        RECT 2054.520 2.400 2054.660 15.650 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1228.730 1670.660 1229.050 1670.720 ;
        RECT 1231.030 1670.660 1231.350 1670.720 ;
        RECT 1228.730 1670.520 1231.350 1670.660 ;
        RECT 1228.730 1670.460 1229.050 1670.520 ;
        RECT 1231.030 1670.460 1231.350 1670.520 ;
        RECT 772.410 1597.560 772.730 1597.620 ;
        RECT 1231.030 1597.560 1231.350 1597.620 ;
        RECT 772.410 1597.420 1231.350 1597.560 ;
        RECT 772.410 1597.360 772.730 1597.420 ;
        RECT 1231.030 1597.360 1231.350 1597.420 ;
      LAYER via ;
        RECT 1228.760 1670.460 1229.020 1670.720 ;
        RECT 1231.060 1670.460 1231.320 1670.720 ;
        RECT 772.440 1597.360 772.700 1597.620 ;
        RECT 1231.060 1597.360 1231.320 1597.620 ;
      LAYER met2 ;
        RECT 1228.660 1700.340 1228.940 1704.000 ;
        RECT 1228.660 1700.000 1228.960 1700.340 ;
        RECT 1228.820 1670.750 1228.960 1700.000 ;
        RECT 1228.760 1670.430 1229.020 1670.750 ;
        RECT 1231.060 1670.430 1231.320 1670.750 ;
        RECT 1231.120 1597.650 1231.260 1670.430 ;
        RECT 772.440 1597.330 772.700 1597.650 ;
        RECT 1231.060 1597.330 1231.320 1597.650 ;
        RECT 772.500 18.090 772.640 1597.330 ;
        RECT 769.740 17.950 772.640 18.090 ;
        RECT 769.740 2.400 769.880 17.950 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1361.670 1678.140 1361.990 1678.200 ;
        RECT 1362.590 1678.140 1362.910 1678.200 ;
        RECT 1361.670 1678.000 1362.910 1678.140 ;
        RECT 1361.670 1677.940 1361.990 1678.000 ;
        RECT 1362.590 1677.940 1362.910 1678.000 ;
        RECT 1361.670 16.220 1361.990 16.280 ;
        RECT 2072.370 16.220 2072.690 16.280 ;
        RECT 1361.670 16.080 2072.690 16.220 ;
        RECT 1361.670 16.020 1361.990 16.080 ;
        RECT 2072.370 16.020 2072.690 16.080 ;
      LAYER via ;
        RECT 1361.700 1677.940 1361.960 1678.200 ;
        RECT 1362.620 1677.940 1362.880 1678.200 ;
        RECT 1361.700 16.020 1361.960 16.280 ;
        RECT 2072.400 16.020 2072.660 16.280 ;
      LAYER met2 ;
        RECT 1362.980 1700.410 1363.260 1704.000 ;
        RECT 1362.680 1700.270 1363.260 1700.410 ;
        RECT 1362.680 1678.230 1362.820 1700.270 ;
        RECT 1362.980 1700.000 1363.260 1700.270 ;
        RECT 1361.700 1677.910 1361.960 1678.230 ;
        RECT 1362.620 1677.910 1362.880 1678.230 ;
        RECT 1361.760 16.310 1361.900 1677.910 ;
        RECT 1361.700 15.990 1361.960 16.310 ;
        RECT 2072.400 15.990 2072.660 16.310 ;
        RECT 2072.460 2.400 2072.600 15.990 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1360.750 1631.900 1361.070 1631.960 ;
        RECT 1364.890 1631.900 1365.210 1631.960 ;
        RECT 1360.750 1631.760 1365.210 1631.900 ;
        RECT 1360.750 1631.700 1361.070 1631.760 ;
        RECT 1364.890 1631.700 1365.210 1631.760 ;
        RECT 1360.750 16.560 1361.070 16.620 ;
        RECT 2089.850 16.560 2090.170 16.620 ;
        RECT 1360.750 16.420 2090.170 16.560 ;
        RECT 1360.750 16.360 1361.070 16.420 ;
        RECT 2089.850 16.360 2090.170 16.420 ;
      LAYER via ;
        RECT 1360.780 1631.700 1361.040 1631.960 ;
        RECT 1364.920 1631.700 1365.180 1631.960 ;
        RECT 1360.780 16.360 1361.040 16.620 ;
        RECT 2089.880 16.360 2090.140 16.620 ;
      LAYER met2 ;
        RECT 1364.820 1700.340 1365.100 1704.000 ;
        RECT 1364.820 1700.000 1365.120 1700.340 ;
        RECT 1364.980 1631.990 1365.120 1700.000 ;
        RECT 1360.780 1631.670 1361.040 1631.990 ;
        RECT 1364.920 1631.670 1365.180 1631.990 ;
        RECT 1360.840 16.650 1360.980 1631.670 ;
        RECT 1360.780 16.330 1361.040 16.650 ;
        RECT 2089.880 16.330 2090.140 16.650 ;
        RECT 2089.940 2.400 2090.080 16.330 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1371.865 1635.485 1372.035 1683.595 ;
        RECT 1371.865 1580.065 1372.035 1628.175 ;
        RECT 1370.945 1187.025 1371.115 1235.135 ;
        RECT 1370.485 607.325 1370.655 655.435 ;
        RECT 1370.485 414.205 1370.655 496.655 ;
        RECT 1371.405 89.845 1371.575 137.955 ;
      LAYER mcon ;
        RECT 1371.865 1683.425 1372.035 1683.595 ;
        RECT 1371.865 1628.005 1372.035 1628.175 ;
        RECT 1370.945 1234.965 1371.115 1235.135 ;
        RECT 1370.485 655.265 1370.655 655.435 ;
        RECT 1370.485 496.485 1370.655 496.655 ;
        RECT 1371.405 137.785 1371.575 137.955 ;
      LAYER met1 ;
        RECT 1366.730 1685.280 1367.050 1685.340 ;
        RECT 1371.790 1685.280 1372.110 1685.340 ;
        RECT 1366.730 1685.140 1372.110 1685.280 ;
        RECT 1366.730 1685.080 1367.050 1685.140 ;
        RECT 1371.790 1685.080 1372.110 1685.140 ;
        RECT 1371.790 1683.580 1372.110 1683.640 ;
        RECT 1371.595 1683.440 1372.110 1683.580 ;
        RECT 1371.790 1683.380 1372.110 1683.440 ;
        RECT 1371.790 1635.640 1372.110 1635.700 ;
        RECT 1371.595 1635.500 1372.110 1635.640 ;
        RECT 1371.790 1635.440 1372.110 1635.500 ;
        RECT 1371.790 1628.160 1372.110 1628.220 ;
        RECT 1371.595 1628.020 1372.110 1628.160 ;
        RECT 1371.790 1627.960 1372.110 1628.020 ;
        RECT 1371.790 1580.220 1372.110 1580.280 ;
        RECT 1371.595 1580.080 1372.110 1580.220 ;
        RECT 1371.790 1580.020 1372.110 1580.080 ;
        RECT 1372.250 1497.940 1372.570 1498.000 ;
        RECT 1371.880 1497.800 1372.570 1497.940 ;
        RECT 1371.880 1497.320 1372.020 1497.800 ;
        RECT 1372.250 1497.740 1372.570 1497.800 ;
        RECT 1371.790 1497.060 1372.110 1497.320 ;
        RECT 1370.870 1249.060 1371.190 1249.120 ;
        RECT 1371.330 1249.060 1371.650 1249.120 ;
        RECT 1370.870 1248.920 1371.650 1249.060 ;
        RECT 1370.870 1248.860 1371.190 1248.920 ;
        RECT 1371.330 1248.860 1371.650 1248.920 ;
        RECT 1370.885 1235.120 1371.175 1235.165 ;
        RECT 1371.330 1235.120 1371.650 1235.180 ;
        RECT 1370.885 1234.980 1371.650 1235.120 ;
        RECT 1370.885 1234.935 1371.175 1234.980 ;
        RECT 1371.330 1234.920 1371.650 1234.980 ;
        RECT 1370.870 1187.180 1371.190 1187.240 ;
        RECT 1370.675 1187.040 1371.190 1187.180 ;
        RECT 1370.870 1186.980 1371.190 1187.040 ;
        RECT 1370.870 1145.160 1371.190 1145.420 ;
        RECT 1370.960 1145.020 1371.100 1145.160 ;
        RECT 1371.790 1145.020 1372.110 1145.080 ;
        RECT 1370.960 1144.880 1372.110 1145.020 ;
        RECT 1371.790 1144.820 1372.110 1144.880 ;
        RECT 1370.870 1069.880 1371.190 1069.940 ;
        RECT 1371.790 1069.880 1372.110 1069.940 ;
        RECT 1370.870 1069.740 1372.110 1069.880 ;
        RECT 1370.870 1069.680 1371.190 1069.740 ;
        RECT 1371.790 1069.680 1372.110 1069.740 ;
        RECT 1370.870 1000.320 1371.190 1000.580 ;
        RECT 1370.960 1000.180 1371.100 1000.320 ;
        RECT 1371.330 1000.180 1371.650 1000.240 ;
        RECT 1370.960 1000.040 1371.650 1000.180 ;
        RECT 1371.330 999.980 1371.650 1000.040 ;
        RECT 1370.870 800.060 1371.190 800.320 ;
        RECT 1370.960 799.640 1371.100 800.060 ;
        RECT 1370.870 799.380 1371.190 799.640 ;
        RECT 1370.425 655.420 1370.715 655.465 ;
        RECT 1370.870 655.420 1371.190 655.480 ;
        RECT 1370.425 655.280 1371.190 655.420 ;
        RECT 1370.425 655.235 1370.715 655.280 ;
        RECT 1370.870 655.220 1371.190 655.280 ;
        RECT 1370.410 607.480 1370.730 607.540 ;
        RECT 1370.215 607.340 1370.730 607.480 ;
        RECT 1370.410 607.280 1370.730 607.340 ;
        RECT 1370.410 559.200 1370.730 559.260 ;
        RECT 1371.330 559.200 1371.650 559.260 ;
        RECT 1370.410 559.060 1371.650 559.200 ;
        RECT 1370.410 559.000 1370.730 559.060 ;
        RECT 1371.330 559.000 1371.650 559.060 ;
        RECT 1370.425 496.640 1370.715 496.685 ;
        RECT 1370.870 496.640 1371.190 496.700 ;
        RECT 1370.425 496.500 1371.190 496.640 ;
        RECT 1370.425 496.455 1370.715 496.500 ;
        RECT 1370.870 496.440 1371.190 496.500 ;
        RECT 1370.425 414.360 1370.715 414.405 ;
        RECT 1370.870 414.360 1371.190 414.420 ;
        RECT 1370.425 414.220 1371.190 414.360 ;
        RECT 1370.425 414.175 1370.715 414.220 ;
        RECT 1370.870 414.160 1371.190 414.220 ;
        RECT 1370.870 383.080 1371.190 383.140 ;
        RECT 1372.250 383.080 1372.570 383.140 ;
        RECT 1370.870 382.940 1372.570 383.080 ;
        RECT 1370.870 382.880 1371.190 382.940 ;
        RECT 1372.250 382.880 1372.570 382.940 ;
        RECT 1371.790 317.800 1372.110 317.860 ;
        RECT 1371.420 317.660 1372.110 317.800 ;
        RECT 1371.420 317.180 1371.560 317.660 ;
        RECT 1371.790 317.600 1372.110 317.660 ;
        RECT 1371.330 316.920 1371.650 317.180 ;
        RECT 1371.330 137.940 1371.650 138.000 ;
        RECT 1371.135 137.800 1371.650 137.940 ;
        RECT 1371.330 137.740 1371.650 137.800 ;
        RECT 1371.330 90.000 1371.650 90.060 ;
        RECT 1371.135 89.860 1371.650 90.000 ;
        RECT 1371.330 89.800 1371.650 89.860 ;
        RECT 1371.330 16.900 1371.650 16.960 ;
        RECT 2107.790 16.900 2108.110 16.960 ;
        RECT 1371.330 16.760 2108.110 16.900 ;
        RECT 1371.330 16.700 1371.650 16.760 ;
        RECT 2107.790 16.700 2108.110 16.760 ;
      LAYER via ;
        RECT 1366.760 1685.080 1367.020 1685.340 ;
        RECT 1371.820 1685.080 1372.080 1685.340 ;
        RECT 1371.820 1683.380 1372.080 1683.640 ;
        RECT 1371.820 1635.440 1372.080 1635.700 ;
        RECT 1371.820 1627.960 1372.080 1628.220 ;
        RECT 1371.820 1580.020 1372.080 1580.280 ;
        RECT 1372.280 1497.740 1372.540 1498.000 ;
        RECT 1371.820 1497.060 1372.080 1497.320 ;
        RECT 1370.900 1248.860 1371.160 1249.120 ;
        RECT 1371.360 1248.860 1371.620 1249.120 ;
        RECT 1371.360 1234.920 1371.620 1235.180 ;
        RECT 1370.900 1186.980 1371.160 1187.240 ;
        RECT 1370.900 1145.160 1371.160 1145.420 ;
        RECT 1371.820 1144.820 1372.080 1145.080 ;
        RECT 1370.900 1069.680 1371.160 1069.940 ;
        RECT 1371.820 1069.680 1372.080 1069.940 ;
        RECT 1370.900 1000.320 1371.160 1000.580 ;
        RECT 1371.360 999.980 1371.620 1000.240 ;
        RECT 1370.900 800.060 1371.160 800.320 ;
        RECT 1370.900 799.380 1371.160 799.640 ;
        RECT 1370.900 655.220 1371.160 655.480 ;
        RECT 1370.440 607.280 1370.700 607.540 ;
        RECT 1370.440 559.000 1370.700 559.260 ;
        RECT 1371.360 559.000 1371.620 559.260 ;
        RECT 1370.900 496.440 1371.160 496.700 ;
        RECT 1370.900 414.160 1371.160 414.420 ;
        RECT 1370.900 382.880 1371.160 383.140 ;
        RECT 1372.280 382.880 1372.540 383.140 ;
        RECT 1371.820 317.600 1372.080 317.860 ;
        RECT 1371.360 316.920 1371.620 317.180 ;
        RECT 1371.360 137.740 1371.620 138.000 ;
        RECT 1371.360 89.800 1371.620 90.060 ;
        RECT 1371.360 16.700 1371.620 16.960 ;
        RECT 2107.820 16.700 2108.080 16.960 ;
      LAYER met2 ;
        RECT 1366.660 1700.340 1366.940 1704.000 ;
        RECT 1366.660 1700.000 1366.960 1700.340 ;
        RECT 1366.820 1685.370 1366.960 1700.000 ;
        RECT 1366.760 1685.050 1367.020 1685.370 ;
        RECT 1371.820 1685.050 1372.080 1685.370 ;
        RECT 1371.880 1683.670 1372.020 1685.050 ;
        RECT 1371.820 1683.350 1372.080 1683.670 ;
        RECT 1371.820 1635.410 1372.080 1635.730 ;
        RECT 1371.880 1628.250 1372.020 1635.410 ;
        RECT 1371.820 1627.930 1372.080 1628.250 ;
        RECT 1371.820 1579.990 1372.080 1580.310 ;
        RECT 1371.880 1556.080 1372.020 1579.990 ;
        RECT 1371.880 1555.940 1372.480 1556.080 ;
        RECT 1372.340 1498.030 1372.480 1555.940 ;
        RECT 1372.280 1497.710 1372.540 1498.030 ;
        RECT 1371.820 1497.030 1372.080 1497.350 ;
        RECT 1371.880 1424.840 1372.020 1497.030 ;
        RECT 1371.420 1424.700 1372.020 1424.840 ;
        RECT 1371.420 1363.130 1371.560 1424.700 ;
        RECT 1370.960 1362.990 1371.560 1363.130 ;
        RECT 1370.960 1249.150 1371.100 1362.990 ;
        RECT 1370.900 1248.830 1371.160 1249.150 ;
        RECT 1371.360 1248.830 1371.620 1249.150 ;
        RECT 1371.420 1235.210 1371.560 1248.830 ;
        RECT 1371.360 1234.890 1371.620 1235.210 ;
        RECT 1370.900 1186.950 1371.160 1187.270 ;
        RECT 1370.960 1145.450 1371.100 1186.950 ;
        RECT 1370.900 1145.130 1371.160 1145.450 ;
        RECT 1371.820 1144.790 1372.080 1145.110 ;
        RECT 1371.880 1069.970 1372.020 1144.790 ;
        RECT 1370.900 1069.650 1371.160 1069.970 ;
        RECT 1371.820 1069.650 1372.080 1069.970 ;
        RECT 1370.960 1000.610 1371.100 1069.650 ;
        RECT 1370.900 1000.290 1371.160 1000.610 ;
        RECT 1371.360 999.950 1371.620 1000.270 ;
        RECT 1371.420 921.130 1371.560 999.950 ;
        RECT 1370.960 920.990 1371.560 921.130 ;
        RECT 1370.960 800.350 1371.100 920.990 ;
        RECT 1370.900 800.030 1371.160 800.350 ;
        RECT 1370.900 799.350 1371.160 799.670 ;
        RECT 1370.960 655.510 1371.100 799.350 ;
        RECT 1370.900 655.190 1371.160 655.510 ;
        RECT 1370.440 607.250 1370.700 607.570 ;
        RECT 1370.500 559.290 1370.640 607.250 ;
        RECT 1370.440 558.970 1370.700 559.290 ;
        RECT 1371.360 558.970 1371.620 559.290 ;
        RECT 1371.420 511.090 1371.560 558.970 ;
        RECT 1370.960 510.950 1371.560 511.090 ;
        RECT 1370.960 496.730 1371.100 510.950 ;
        RECT 1370.900 496.410 1371.160 496.730 ;
        RECT 1370.900 414.130 1371.160 414.450 ;
        RECT 1370.960 383.170 1371.100 414.130 ;
        RECT 1370.900 382.850 1371.160 383.170 ;
        RECT 1372.280 382.850 1372.540 383.170 ;
        RECT 1372.340 358.770 1372.480 382.850 ;
        RECT 1371.880 358.630 1372.480 358.770 ;
        RECT 1371.880 317.890 1372.020 358.630 ;
        RECT 1371.820 317.570 1372.080 317.890 ;
        RECT 1371.360 316.890 1371.620 317.210 ;
        RECT 1371.420 138.030 1371.560 316.890 ;
        RECT 1371.360 137.710 1371.620 138.030 ;
        RECT 1371.360 89.770 1371.620 90.090 ;
        RECT 1371.420 16.990 1371.560 89.770 ;
        RECT 1371.360 16.670 1371.620 16.990 ;
        RECT 2107.820 16.670 2108.080 16.990 ;
        RECT 2107.880 2.400 2108.020 16.670 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1369.105 903.805 1369.275 921.315 ;
        RECT 1369.565 552.245 1369.735 600.355 ;
        RECT 1369.565 317.645 1369.735 383.095 ;
      LAYER mcon ;
        RECT 1369.105 921.145 1369.275 921.315 ;
        RECT 1369.565 600.185 1369.735 600.355 ;
        RECT 1369.565 382.925 1369.735 383.095 ;
      LAYER met1 ;
        RECT 1369.030 1448.980 1369.350 1449.040 ;
        RECT 1369.490 1448.980 1369.810 1449.040 ;
        RECT 1369.030 1448.840 1369.810 1448.980 ;
        RECT 1369.030 1448.780 1369.350 1448.840 ;
        RECT 1369.490 1448.780 1369.810 1448.840 ;
        RECT 1369.490 1014.460 1369.810 1014.520 ;
        RECT 1369.950 1014.460 1370.270 1014.520 ;
        RECT 1369.490 1014.320 1370.270 1014.460 ;
        RECT 1369.490 1014.260 1369.810 1014.320 ;
        RECT 1369.950 1014.260 1370.270 1014.320 ;
        RECT 1369.045 921.300 1369.335 921.345 ;
        RECT 1369.490 921.300 1369.810 921.360 ;
        RECT 1369.045 921.160 1369.810 921.300 ;
        RECT 1369.045 921.115 1369.335 921.160 ;
        RECT 1369.490 921.100 1369.810 921.160 ;
        RECT 1369.030 903.960 1369.350 904.020 ;
        RECT 1368.835 903.820 1369.350 903.960 ;
        RECT 1369.030 903.760 1369.350 903.820 ;
        RECT 1369.030 855.340 1369.350 855.400 ;
        RECT 1369.490 855.340 1369.810 855.400 ;
        RECT 1369.030 855.200 1369.810 855.340 ;
        RECT 1369.030 855.140 1369.350 855.200 ;
        RECT 1369.490 855.140 1369.810 855.200 ;
        RECT 1369.030 710.840 1369.350 710.900 ;
        RECT 1369.490 710.840 1369.810 710.900 ;
        RECT 1369.030 710.700 1369.810 710.840 ;
        RECT 1369.030 710.640 1369.350 710.700 ;
        RECT 1369.490 710.640 1369.810 710.700 ;
        RECT 1369.030 669.360 1369.350 669.420 ;
        RECT 1369.950 669.360 1370.270 669.420 ;
        RECT 1369.030 669.220 1370.270 669.360 ;
        RECT 1369.030 669.160 1369.350 669.220 ;
        RECT 1369.950 669.160 1370.270 669.220 ;
        RECT 1369.490 600.340 1369.810 600.400 ;
        RECT 1369.295 600.200 1369.810 600.340 ;
        RECT 1369.490 600.140 1369.810 600.200 ;
        RECT 1369.505 552.400 1369.795 552.445 ;
        RECT 1369.950 552.400 1370.270 552.460 ;
        RECT 1369.505 552.260 1370.270 552.400 ;
        RECT 1369.505 552.215 1369.795 552.260 ;
        RECT 1369.950 552.200 1370.270 552.260 ;
        RECT 1369.030 462.300 1369.350 462.360 ;
        RECT 1369.950 462.300 1370.270 462.360 ;
        RECT 1369.030 462.160 1370.270 462.300 ;
        RECT 1369.030 462.100 1369.350 462.160 ;
        RECT 1369.950 462.100 1370.270 462.160 ;
        RECT 1369.505 383.080 1369.795 383.125 ;
        RECT 1370.410 383.080 1370.730 383.140 ;
        RECT 1369.505 382.940 1370.730 383.080 ;
        RECT 1369.505 382.895 1369.795 382.940 ;
        RECT 1370.410 382.880 1370.730 382.940 ;
        RECT 1369.490 317.800 1369.810 317.860 ;
        RECT 1369.295 317.660 1369.810 317.800 ;
        RECT 1369.490 317.600 1369.810 317.660 ;
        RECT 1369.490 241.640 1369.810 241.700 ;
        RECT 1369.950 241.640 1370.270 241.700 ;
        RECT 1369.490 241.500 1370.270 241.640 ;
        RECT 1369.490 241.440 1369.810 241.500 ;
        RECT 1369.950 241.440 1370.270 241.500 ;
        RECT 1369.030 20.640 1369.350 20.700 ;
        RECT 2125.270 20.640 2125.590 20.700 ;
        RECT 1369.030 20.500 2125.590 20.640 ;
        RECT 1369.030 20.440 1369.350 20.500 ;
        RECT 2125.270 20.440 2125.590 20.500 ;
      LAYER via ;
        RECT 1369.060 1448.780 1369.320 1449.040 ;
        RECT 1369.520 1448.780 1369.780 1449.040 ;
        RECT 1369.520 1014.260 1369.780 1014.520 ;
        RECT 1369.980 1014.260 1370.240 1014.520 ;
        RECT 1369.520 921.100 1369.780 921.360 ;
        RECT 1369.060 903.760 1369.320 904.020 ;
        RECT 1369.060 855.140 1369.320 855.400 ;
        RECT 1369.520 855.140 1369.780 855.400 ;
        RECT 1369.060 710.640 1369.320 710.900 ;
        RECT 1369.520 710.640 1369.780 710.900 ;
        RECT 1369.060 669.160 1369.320 669.420 ;
        RECT 1369.980 669.160 1370.240 669.420 ;
        RECT 1369.520 600.140 1369.780 600.400 ;
        RECT 1369.980 552.200 1370.240 552.460 ;
        RECT 1369.060 462.100 1369.320 462.360 ;
        RECT 1369.980 462.100 1370.240 462.360 ;
        RECT 1370.440 382.880 1370.700 383.140 ;
        RECT 1369.520 317.600 1369.780 317.860 ;
        RECT 1369.520 241.440 1369.780 241.700 ;
        RECT 1369.980 241.440 1370.240 241.700 ;
        RECT 1369.060 20.440 1369.320 20.700 ;
        RECT 2125.300 20.440 2125.560 20.700 ;
      LAYER met2 ;
        RECT 1368.500 1700.410 1368.780 1704.000 ;
        RECT 1368.200 1700.270 1368.780 1700.410 ;
        RECT 1368.200 1684.885 1368.340 1700.270 ;
        RECT 1368.500 1700.000 1368.780 1700.270 ;
        RECT 1368.130 1684.515 1368.410 1684.885 ;
        RECT 1369.050 1683.835 1369.330 1684.205 ;
        RECT 1369.120 1449.070 1369.260 1683.835 ;
        RECT 1369.060 1448.750 1369.320 1449.070 ;
        RECT 1369.520 1448.750 1369.780 1449.070 ;
        RECT 1369.580 1072.770 1369.720 1448.750 ;
        RECT 1369.580 1072.630 1370.180 1072.770 ;
        RECT 1370.040 1014.550 1370.180 1072.630 ;
        RECT 1369.520 1014.230 1369.780 1014.550 ;
        RECT 1369.980 1014.230 1370.240 1014.550 ;
        RECT 1369.580 921.390 1369.720 1014.230 ;
        RECT 1369.520 921.070 1369.780 921.390 ;
        RECT 1369.060 903.730 1369.320 904.050 ;
        RECT 1369.120 855.430 1369.260 903.730 ;
        RECT 1369.060 855.110 1369.320 855.430 ;
        RECT 1369.520 855.110 1369.780 855.430 ;
        RECT 1369.580 710.930 1369.720 855.110 ;
        RECT 1369.060 710.610 1369.320 710.930 ;
        RECT 1369.520 710.610 1369.780 710.930 ;
        RECT 1369.120 669.450 1369.260 710.610 ;
        RECT 1369.060 669.130 1369.320 669.450 ;
        RECT 1369.980 669.130 1370.240 669.450 ;
        RECT 1370.040 644.370 1370.180 669.130 ;
        RECT 1369.580 644.230 1370.180 644.370 ;
        RECT 1369.580 600.430 1369.720 644.230 ;
        RECT 1369.520 600.110 1369.780 600.430 ;
        RECT 1369.980 552.170 1370.240 552.490 ;
        RECT 1370.040 462.390 1370.180 552.170 ;
        RECT 1369.060 462.070 1369.320 462.390 ;
        RECT 1369.980 462.070 1370.240 462.390 ;
        RECT 1369.120 455.445 1369.260 462.070 ;
        RECT 1369.050 455.075 1369.330 455.445 ;
        RECT 1370.430 455.075 1370.710 455.445 ;
        RECT 1370.500 383.170 1370.640 455.075 ;
        RECT 1370.440 382.850 1370.700 383.170 ;
        RECT 1369.520 317.570 1369.780 317.890 ;
        RECT 1369.580 317.290 1369.720 317.570 ;
        RECT 1369.580 317.150 1370.180 317.290 ;
        RECT 1370.040 241.730 1370.180 317.150 ;
        RECT 1369.520 241.410 1369.780 241.730 ;
        RECT 1369.980 241.410 1370.240 241.730 ;
        RECT 1369.580 169.050 1369.720 241.410 ;
        RECT 1369.120 168.910 1369.720 169.050 ;
        RECT 1369.120 20.730 1369.260 168.910 ;
        RECT 1369.060 20.410 1369.320 20.730 ;
        RECT 2125.300 20.410 2125.560 20.730 ;
        RECT 2125.360 14.010 2125.500 20.410 ;
        RECT 2125.360 13.870 2125.960 14.010 ;
        RECT 2125.820 2.400 2125.960 13.870 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
      LAYER via2 ;
        RECT 1368.130 1684.560 1368.410 1684.840 ;
        RECT 1369.050 1683.880 1369.330 1684.160 ;
        RECT 1369.050 455.120 1369.330 455.400 ;
        RECT 1370.430 455.120 1370.710 455.400 ;
      LAYER met3 ;
        RECT 1368.105 1684.850 1368.435 1684.865 ;
        RECT 1368.105 1684.535 1368.650 1684.850 ;
        RECT 1368.350 1684.170 1368.650 1684.535 ;
        RECT 1369.025 1684.170 1369.355 1684.185 ;
        RECT 1368.350 1683.870 1369.355 1684.170 ;
        RECT 1369.025 1683.855 1369.355 1683.870 ;
        RECT 1369.025 455.410 1369.355 455.425 ;
        RECT 1370.405 455.410 1370.735 455.425 ;
        RECT 1369.025 455.110 1370.735 455.410 ;
        RECT 1369.025 455.095 1369.355 455.110 ;
        RECT 1370.405 455.095 1370.735 455.110 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1368.185 1483.505 1368.355 1545.555 ;
      LAYER mcon ;
        RECT 1368.185 1545.385 1368.355 1545.555 ;
      LAYER met1 ;
        RECT 1368.110 1556.080 1368.430 1556.140 ;
        RECT 1369.950 1556.080 1370.270 1556.140 ;
        RECT 1368.110 1555.940 1370.270 1556.080 ;
        RECT 1368.110 1555.880 1368.430 1555.940 ;
        RECT 1369.950 1555.880 1370.270 1555.940 ;
        RECT 1368.110 1545.540 1368.430 1545.600 ;
        RECT 1367.915 1545.400 1368.430 1545.540 ;
        RECT 1368.110 1545.340 1368.430 1545.400 ;
        RECT 1368.110 1483.660 1368.430 1483.720 ;
        RECT 1367.915 1483.520 1368.430 1483.660 ;
        RECT 1368.110 1483.460 1368.430 1483.520 ;
        RECT 1368.110 1317.880 1368.430 1318.140 ;
        RECT 1368.200 1317.740 1368.340 1317.880 ;
        RECT 1368.570 1317.740 1368.890 1317.800 ;
        RECT 1368.200 1317.600 1368.890 1317.740 ;
        RECT 1368.570 1317.540 1368.890 1317.600 ;
        RECT 1368.570 1256.000 1368.890 1256.260 ;
        RECT 1368.660 1255.520 1368.800 1256.000 ;
        RECT 1369.030 1255.520 1369.350 1255.580 ;
        RECT 1368.660 1255.380 1369.350 1255.520 ;
        RECT 1369.030 1255.320 1369.350 1255.380 ;
        RECT 1368.570 1207.580 1368.890 1207.640 ;
        RECT 1369.030 1207.580 1369.350 1207.640 ;
        RECT 1368.570 1207.440 1369.350 1207.580 ;
        RECT 1368.570 1207.380 1368.890 1207.440 ;
        RECT 1369.030 1207.380 1369.350 1207.440 ;
        RECT 1368.570 917.900 1368.890 917.960 ;
        RECT 1369.030 917.900 1369.350 917.960 ;
        RECT 1368.570 917.760 1369.350 917.900 ;
        RECT 1368.570 917.700 1368.890 917.760 ;
        RECT 1369.030 917.700 1369.350 917.760 ;
        RECT 1368.110 821.140 1368.430 821.400 ;
        RECT 1368.200 820.660 1368.340 821.140 ;
        RECT 1368.570 820.660 1368.890 820.720 ;
        RECT 1368.200 820.520 1368.890 820.660 ;
        RECT 1368.570 820.460 1368.890 820.520 ;
        RECT 1368.110 710.840 1368.430 710.900 ;
        RECT 1368.570 710.840 1368.890 710.900 ;
        RECT 1368.110 710.700 1368.890 710.840 ;
        RECT 1368.110 710.640 1368.430 710.700 ;
        RECT 1368.570 710.640 1368.890 710.700 ;
        RECT 1368.110 372.880 1368.430 372.940 ;
        RECT 1368.570 372.880 1368.890 372.940 ;
        RECT 1368.110 372.740 1368.890 372.880 ;
        RECT 1368.110 372.680 1368.430 372.740 ;
        RECT 1368.570 372.680 1368.890 372.740 ;
        RECT 1368.110 331.540 1368.430 331.800 ;
        RECT 1368.200 331.120 1368.340 331.540 ;
        RECT 1368.110 330.860 1368.430 331.120 ;
        RECT 1368.110 293.320 1368.430 293.380 ;
        RECT 1369.490 293.320 1369.810 293.380 ;
        RECT 1368.110 293.180 1369.810 293.320 ;
        RECT 1368.110 293.120 1368.430 293.180 ;
        RECT 1369.490 293.120 1369.810 293.180 ;
        RECT 1368.110 186.220 1368.430 186.280 ;
        RECT 1368.570 186.220 1368.890 186.280 ;
        RECT 1368.110 186.080 1368.890 186.220 ;
        RECT 1368.110 186.020 1368.430 186.080 ;
        RECT 1368.570 186.020 1368.890 186.080 ;
        RECT 1368.110 20.300 1368.430 20.360 ;
        RECT 2143.670 20.300 2143.990 20.360 ;
        RECT 1368.110 20.160 2143.990 20.300 ;
        RECT 1368.110 20.100 1368.430 20.160 ;
        RECT 2143.670 20.100 2143.990 20.160 ;
      LAYER via ;
        RECT 1368.140 1555.880 1368.400 1556.140 ;
        RECT 1369.980 1555.880 1370.240 1556.140 ;
        RECT 1368.140 1545.340 1368.400 1545.600 ;
        RECT 1368.140 1483.460 1368.400 1483.720 ;
        RECT 1368.140 1317.880 1368.400 1318.140 ;
        RECT 1368.600 1317.540 1368.860 1317.800 ;
        RECT 1368.600 1256.000 1368.860 1256.260 ;
        RECT 1369.060 1255.320 1369.320 1255.580 ;
        RECT 1368.600 1207.380 1368.860 1207.640 ;
        RECT 1369.060 1207.380 1369.320 1207.640 ;
        RECT 1368.600 917.700 1368.860 917.960 ;
        RECT 1369.060 917.700 1369.320 917.960 ;
        RECT 1368.140 821.140 1368.400 821.400 ;
        RECT 1368.600 820.460 1368.860 820.720 ;
        RECT 1368.140 710.640 1368.400 710.900 ;
        RECT 1368.600 710.640 1368.860 710.900 ;
        RECT 1368.140 372.680 1368.400 372.940 ;
        RECT 1368.600 372.680 1368.860 372.940 ;
        RECT 1368.140 331.540 1368.400 331.800 ;
        RECT 1368.140 330.860 1368.400 331.120 ;
        RECT 1368.140 293.120 1368.400 293.380 ;
        RECT 1369.520 293.120 1369.780 293.380 ;
        RECT 1368.140 186.020 1368.400 186.280 ;
        RECT 1368.600 186.020 1368.860 186.280 ;
        RECT 1368.140 20.100 1368.400 20.360 ;
        RECT 2143.700 20.100 2143.960 20.360 ;
      LAYER met2 ;
        RECT 1370.340 1700.410 1370.620 1704.000 ;
        RECT 1370.040 1700.270 1370.620 1700.410 ;
        RECT 1370.040 1556.170 1370.180 1700.270 ;
        RECT 1370.340 1700.000 1370.620 1700.270 ;
        RECT 1368.140 1555.850 1368.400 1556.170 ;
        RECT 1369.980 1555.850 1370.240 1556.170 ;
        RECT 1368.200 1545.630 1368.340 1555.850 ;
        RECT 1368.140 1545.310 1368.400 1545.630 ;
        RECT 1368.140 1483.430 1368.400 1483.750 ;
        RECT 1368.200 1318.170 1368.340 1483.430 ;
        RECT 1368.140 1317.850 1368.400 1318.170 ;
        RECT 1368.600 1317.510 1368.860 1317.830 ;
        RECT 1368.660 1256.290 1368.800 1317.510 ;
        RECT 1368.600 1255.970 1368.860 1256.290 ;
        RECT 1369.060 1255.290 1369.320 1255.610 ;
        RECT 1369.120 1207.670 1369.260 1255.290 ;
        RECT 1368.600 1207.350 1368.860 1207.670 ;
        RECT 1369.060 1207.350 1369.320 1207.670 ;
        RECT 1368.660 976.210 1368.800 1207.350 ;
        RECT 1368.660 976.070 1369.260 976.210 ;
        RECT 1369.120 917.990 1369.260 976.070 ;
        RECT 1368.600 917.670 1368.860 917.990 ;
        RECT 1369.060 917.670 1369.320 917.990 ;
        RECT 1368.660 879.650 1368.800 917.670 ;
        RECT 1368.200 879.510 1368.800 879.650 ;
        RECT 1368.200 821.430 1368.340 879.510 ;
        RECT 1368.140 821.110 1368.400 821.430 ;
        RECT 1368.600 820.430 1368.860 820.750 ;
        RECT 1368.660 710.930 1368.800 820.430 ;
        RECT 1368.140 710.610 1368.400 710.930 ;
        RECT 1368.600 710.610 1368.860 710.930 ;
        RECT 1368.200 559.370 1368.340 710.610 ;
        RECT 1368.200 559.230 1368.800 559.370 ;
        RECT 1368.660 372.970 1368.800 559.230 ;
        RECT 1368.140 372.650 1368.400 372.970 ;
        RECT 1368.600 372.650 1368.860 372.970 ;
        RECT 1368.200 331.830 1368.340 372.650 ;
        RECT 1368.140 331.510 1368.400 331.830 ;
        RECT 1368.140 330.830 1368.400 331.150 ;
        RECT 1368.200 293.410 1368.340 330.830 ;
        RECT 1368.140 293.090 1368.400 293.410 ;
        RECT 1369.520 293.090 1369.780 293.410 ;
        RECT 1369.580 252.010 1369.720 293.090 ;
        RECT 1369.120 251.870 1369.720 252.010 ;
        RECT 1369.120 241.810 1369.260 251.870 ;
        RECT 1368.660 241.670 1369.260 241.810 ;
        RECT 1368.660 186.310 1368.800 241.670 ;
        RECT 1368.140 185.990 1368.400 186.310 ;
        RECT 1368.600 185.990 1368.860 186.310 ;
        RECT 1368.200 20.390 1368.340 185.990 ;
        RECT 1368.140 20.070 1368.400 20.390 ;
        RECT 2143.700 20.070 2143.960 20.390 ;
        RECT 2143.760 2.400 2143.900 20.070 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1372.250 1683.920 1372.570 1683.980 ;
        RECT 1370.040 1683.780 1372.570 1683.920 ;
        RECT 1367.650 1683.580 1367.970 1683.640 ;
        RECT 1370.040 1683.580 1370.180 1683.780 ;
        RECT 1372.250 1683.720 1372.570 1683.780 ;
        RECT 1367.650 1683.440 1370.180 1683.580 ;
        RECT 1367.650 1683.380 1367.970 1683.440 ;
        RECT 1367.650 19.960 1367.970 20.020 ;
        RECT 2161.610 19.960 2161.930 20.020 ;
        RECT 1367.650 19.820 2161.930 19.960 ;
        RECT 1367.650 19.760 1367.970 19.820 ;
        RECT 2161.610 19.760 2161.930 19.820 ;
      LAYER via ;
        RECT 1367.680 1683.380 1367.940 1683.640 ;
        RECT 1372.280 1683.720 1372.540 1683.980 ;
        RECT 1367.680 19.760 1367.940 20.020 ;
        RECT 2161.640 19.760 2161.900 20.020 ;
      LAYER met2 ;
        RECT 1372.180 1700.340 1372.460 1704.000 ;
        RECT 1372.180 1700.000 1372.480 1700.340 ;
        RECT 1372.340 1684.010 1372.480 1700.000 ;
        RECT 1372.280 1683.690 1372.540 1684.010 ;
        RECT 1367.680 1683.350 1367.940 1683.670 ;
        RECT 1367.740 20.050 1367.880 1683.350 ;
        RECT 1367.680 19.730 1367.940 20.050 ;
        RECT 2161.640 19.730 2161.900 20.050 ;
        RECT 2161.700 2.400 2161.840 19.730 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1374.090 1665.220 1374.410 1665.280 ;
        RECT 1378.690 1665.220 1379.010 1665.280 ;
        RECT 1374.090 1665.080 1379.010 1665.220 ;
        RECT 1374.090 1665.020 1374.410 1665.080 ;
        RECT 1378.690 1665.020 1379.010 1665.080 ;
        RECT 1378.690 19.620 1379.010 19.680 ;
        RECT 2179.090 19.620 2179.410 19.680 ;
        RECT 1378.690 19.480 2179.410 19.620 ;
        RECT 1378.690 19.420 1379.010 19.480 ;
        RECT 2179.090 19.420 2179.410 19.480 ;
      LAYER via ;
        RECT 1374.120 1665.020 1374.380 1665.280 ;
        RECT 1378.720 1665.020 1378.980 1665.280 ;
        RECT 1378.720 19.420 1378.980 19.680 ;
        RECT 2179.120 19.420 2179.380 19.680 ;
      LAYER met2 ;
        RECT 1374.020 1700.340 1374.300 1704.000 ;
        RECT 1374.020 1700.000 1374.320 1700.340 ;
        RECT 1374.180 1665.310 1374.320 1700.000 ;
        RECT 1374.120 1664.990 1374.380 1665.310 ;
        RECT 1378.720 1664.990 1378.980 1665.310 ;
        RECT 1378.780 19.710 1378.920 1664.990 ;
        RECT 1378.720 19.390 1378.980 19.710 ;
        RECT 2179.120 19.390 2179.380 19.710 ;
        RECT 2179.180 2.400 2179.320 19.390 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1375.470 19.280 1375.790 19.340 ;
        RECT 2197.030 19.280 2197.350 19.340 ;
        RECT 1375.470 19.140 2197.350 19.280 ;
        RECT 1375.470 19.080 1375.790 19.140 ;
        RECT 2197.030 19.080 2197.350 19.140 ;
      LAYER via ;
        RECT 1375.500 19.080 1375.760 19.340 ;
        RECT 2197.060 19.080 2197.320 19.340 ;
      LAYER met2 ;
        RECT 1375.400 1700.340 1375.680 1704.000 ;
        RECT 1375.400 1700.000 1375.700 1700.340 ;
        RECT 1375.560 19.370 1375.700 1700.000 ;
        RECT 1375.500 19.050 1375.760 19.370 ;
        RECT 2197.060 19.050 2197.320 19.370 ;
        RECT 2197.120 2.400 2197.260 19.050 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1376.390 1683.920 1376.710 1683.980 ;
        RECT 1377.310 1683.920 1377.630 1683.980 ;
        RECT 1376.390 1683.780 1377.630 1683.920 ;
        RECT 1376.390 1683.720 1376.710 1683.780 ;
        RECT 1377.310 1683.720 1377.630 1683.780 ;
        RECT 1376.850 18.940 1377.170 19.000 ;
        RECT 2214.970 18.940 2215.290 19.000 ;
        RECT 1376.850 18.800 2215.290 18.940 ;
        RECT 1376.850 18.740 1377.170 18.800 ;
        RECT 2214.970 18.740 2215.290 18.800 ;
      LAYER via ;
        RECT 1376.420 1683.720 1376.680 1683.980 ;
        RECT 1377.340 1683.720 1377.600 1683.980 ;
        RECT 1376.880 18.740 1377.140 19.000 ;
        RECT 2215.000 18.740 2215.260 19.000 ;
      LAYER met2 ;
        RECT 1377.240 1700.340 1377.520 1704.000 ;
        RECT 1377.240 1700.000 1377.540 1700.340 ;
        RECT 1377.400 1684.010 1377.540 1700.000 ;
        RECT 1376.420 1683.690 1376.680 1684.010 ;
        RECT 1377.340 1683.690 1377.600 1684.010 ;
        RECT 1376.480 41.890 1376.620 1683.690 ;
        RECT 1376.480 41.750 1377.080 41.890 ;
        RECT 1376.940 19.030 1377.080 41.750 ;
        RECT 1376.880 18.710 1377.140 19.030 ;
        RECT 2215.000 18.710 2215.260 19.030 ;
        RECT 2215.060 2.400 2215.200 18.710 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1379.150 1656.720 1379.470 1656.780 ;
        RECT 1375.100 1656.580 1379.470 1656.720 ;
        RECT 1375.100 1656.100 1375.240 1656.580 ;
        RECT 1379.150 1656.520 1379.470 1656.580 ;
        RECT 1375.010 1655.840 1375.330 1656.100 ;
        RECT 1375.010 18.600 1375.330 18.660 ;
        RECT 2232.910 18.600 2233.230 18.660 ;
        RECT 1375.010 18.460 2233.230 18.600 ;
        RECT 1375.010 18.400 1375.330 18.460 ;
        RECT 2232.910 18.400 2233.230 18.460 ;
      LAYER via ;
        RECT 1379.180 1656.520 1379.440 1656.780 ;
        RECT 1375.040 1655.840 1375.300 1656.100 ;
        RECT 1375.040 18.400 1375.300 18.660 ;
        RECT 2232.940 18.400 2233.200 18.660 ;
      LAYER met2 ;
        RECT 1379.080 1700.340 1379.360 1704.000 ;
        RECT 1379.080 1700.000 1379.380 1700.340 ;
        RECT 1379.240 1656.810 1379.380 1700.000 ;
        RECT 1379.180 1656.490 1379.440 1656.810 ;
        RECT 1375.040 1655.810 1375.300 1656.130 ;
        RECT 1375.100 18.690 1375.240 1655.810 ;
        RECT 1375.040 18.370 1375.300 18.690 ;
        RECT 2232.940 18.370 2233.200 18.690 ;
        RECT 2233.000 2.400 2233.140 18.370 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.110 1563.220 793.430 1563.280 ;
        RECT 1230.570 1563.220 1230.890 1563.280 ;
        RECT 793.110 1563.080 1230.890 1563.220 ;
        RECT 793.110 1563.020 793.430 1563.080 ;
        RECT 1230.570 1563.020 1230.890 1563.080 ;
      LAYER via ;
        RECT 793.140 1563.020 793.400 1563.280 ;
        RECT 1230.600 1563.020 1230.860 1563.280 ;
      LAYER met2 ;
        RECT 1230.500 1700.340 1230.780 1704.000 ;
        RECT 1230.500 1700.000 1230.800 1700.340 ;
        RECT 1230.660 1563.310 1230.800 1700.000 ;
        RECT 793.140 1562.990 793.400 1563.310 ;
        RECT 1230.600 1562.990 1230.860 1563.310 ;
        RECT 793.200 18.090 793.340 1562.990 ;
        RECT 787.680 17.950 793.340 18.090 ;
        RECT 787.680 2.400 787.820 17.950 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1381.450 1670.660 1381.770 1670.720 ;
        RECT 1382.370 1670.660 1382.690 1670.720 ;
        RECT 1381.450 1670.520 1382.690 1670.660 ;
        RECT 1381.450 1670.460 1381.770 1670.520 ;
        RECT 1382.370 1670.460 1382.690 1670.520 ;
        RECT 1382.830 18.260 1383.150 18.320 ;
        RECT 2250.850 18.260 2251.170 18.320 ;
        RECT 1382.830 18.120 2251.170 18.260 ;
        RECT 1382.830 18.060 1383.150 18.120 ;
        RECT 2250.850 18.060 2251.170 18.120 ;
      LAYER via ;
        RECT 1381.480 1670.460 1381.740 1670.720 ;
        RECT 1382.400 1670.460 1382.660 1670.720 ;
        RECT 1382.860 18.060 1383.120 18.320 ;
        RECT 2250.880 18.060 2251.140 18.320 ;
      LAYER met2 ;
        RECT 1380.920 1700.410 1381.200 1704.000 ;
        RECT 1380.920 1700.270 1381.680 1700.410 ;
        RECT 1380.920 1700.000 1381.200 1700.270 ;
        RECT 1381.540 1670.750 1381.680 1700.270 ;
        RECT 1381.480 1670.430 1381.740 1670.750 ;
        RECT 1382.400 1670.430 1382.660 1670.750 ;
        RECT 1382.460 40.530 1382.600 1670.430 ;
        RECT 1382.460 40.390 1383.060 40.530 ;
        RECT 1382.920 18.350 1383.060 40.390 ;
        RECT 1382.860 18.030 1383.120 18.350 ;
        RECT 2250.880 18.030 2251.140 18.350 ;
        RECT 2250.940 2.400 2251.080 18.030 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1381.910 17.920 1382.230 17.980 ;
        RECT 2268.330 17.920 2268.650 17.980 ;
        RECT 1381.910 17.780 2268.650 17.920 ;
        RECT 1381.910 17.720 1382.230 17.780 ;
        RECT 2268.330 17.720 2268.650 17.780 ;
      LAYER via ;
        RECT 1381.940 17.720 1382.200 17.980 ;
        RECT 2268.360 17.720 2268.620 17.980 ;
      LAYER met2 ;
        RECT 1382.760 1700.340 1383.040 1704.000 ;
        RECT 1382.760 1700.000 1383.060 1700.340 ;
        RECT 1382.920 1671.170 1383.060 1700.000 ;
        RECT 1382.000 1671.030 1383.060 1671.170 ;
        RECT 1382.000 18.010 1382.140 1671.030 ;
        RECT 1381.940 17.690 1382.200 18.010 ;
        RECT 2268.360 17.690 2268.620 18.010 ;
        RECT 2268.420 2.400 2268.560 17.690 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1385.205 1676.965 1385.375 1692.775 ;
        RECT 1386.125 1324.725 1386.295 1373.175 ;
        RECT 1386.125 1234.965 1386.295 1276.275 ;
        RECT 1386.125 1187.025 1386.295 1207.595 ;
        RECT 1385.665 938.485 1385.835 986.595 ;
        RECT 1385.665 697.085 1385.835 745.195 ;
        RECT 1386.125 511.105 1386.295 579.955 ;
        RECT 1385.665 372.725 1385.835 420.835 ;
        RECT 1385.665 317.645 1385.835 365.415 ;
      LAYER mcon ;
        RECT 1385.205 1692.605 1385.375 1692.775 ;
        RECT 1386.125 1373.005 1386.295 1373.175 ;
        RECT 1386.125 1276.105 1386.295 1276.275 ;
        RECT 1386.125 1207.425 1386.295 1207.595 ;
        RECT 1385.665 986.425 1385.835 986.595 ;
        RECT 1385.665 745.025 1385.835 745.195 ;
        RECT 1386.125 579.785 1386.295 579.955 ;
        RECT 1385.665 420.665 1385.835 420.835 ;
        RECT 1385.665 365.245 1385.835 365.415 ;
      LAYER met1 ;
        RECT 1385.130 1692.760 1385.450 1692.820 ;
        RECT 1384.935 1692.620 1385.450 1692.760 ;
        RECT 1385.130 1692.560 1385.450 1692.620 ;
        RECT 1385.130 1677.120 1385.450 1677.180 ;
        RECT 1384.935 1676.980 1385.450 1677.120 ;
        RECT 1385.130 1676.920 1385.450 1676.980 ;
        RECT 1385.130 1635.300 1385.450 1635.360 ;
        RECT 1385.590 1635.300 1385.910 1635.360 ;
        RECT 1385.130 1635.160 1385.910 1635.300 ;
        RECT 1385.130 1635.100 1385.450 1635.160 ;
        RECT 1385.590 1635.100 1385.910 1635.160 ;
        RECT 1385.590 1452.380 1385.910 1452.440 ;
        RECT 1386.510 1452.380 1386.830 1452.440 ;
        RECT 1385.590 1452.240 1386.830 1452.380 ;
        RECT 1385.590 1452.180 1385.910 1452.240 ;
        RECT 1386.510 1452.180 1386.830 1452.240 ;
        RECT 1385.590 1448.980 1385.910 1449.040 ;
        RECT 1386.510 1448.980 1386.830 1449.040 ;
        RECT 1385.590 1448.840 1386.830 1448.980 ;
        RECT 1385.590 1448.780 1385.910 1448.840 ;
        RECT 1386.510 1448.780 1386.830 1448.840 ;
        RECT 1386.050 1373.160 1386.370 1373.220 ;
        RECT 1385.855 1373.020 1386.370 1373.160 ;
        RECT 1386.050 1372.960 1386.370 1373.020 ;
        RECT 1386.050 1324.880 1386.370 1324.940 ;
        RECT 1385.855 1324.740 1386.370 1324.880 ;
        RECT 1386.050 1324.680 1386.370 1324.740 ;
        RECT 1386.050 1276.260 1386.370 1276.320 ;
        RECT 1385.855 1276.120 1386.370 1276.260 ;
        RECT 1386.050 1276.060 1386.370 1276.120 ;
        RECT 1386.050 1235.120 1386.370 1235.180 ;
        RECT 1385.855 1234.980 1386.370 1235.120 ;
        RECT 1386.050 1234.920 1386.370 1234.980 ;
        RECT 1386.050 1207.580 1386.370 1207.640 ;
        RECT 1385.855 1207.440 1386.370 1207.580 ;
        RECT 1386.050 1207.380 1386.370 1207.440 ;
        RECT 1386.050 1187.180 1386.370 1187.240 ;
        RECT 1385.855 1187.040 1386.370 1187.180 ;
        RECT 1386.050 1186.980 1386.370 1187.040 ;
        RECT 1385.590 1048.800 1385.910 1048.860 ;
        RECT 1386.050 1048.800 1386.370 1048.860 ;
        RECT 1385.590 1048.660 1386.370 1048.800 ;
        RECT 1385.590 1048.600 1385.910 1048.660 ;
        RECT 1386.050 1048.600 1386.370 1048.660 ;
        RECT 1385.590 1041.660 1385.910 1041.720 ;
        RECT 1386.050 1041.660 1386.370 1041.720 ;
        RECT 1385.590 1041.520 1386.370 1041.660 ;
        RECT 1385.590 1041.460 1385.910 1041.520 ;
        RECT 1386.050 1041.460 1386.370 1041.520 ;
        RECT 1385.590 986.580 1385.910 986.640 ;
        RECT 1385.395 986.440 1385.910 986.580 ;
        RECT 1385.590 986.380 1385.910 986.440 ;
        RECT 1385.590 938.640 1385.910 938.700 ;
        RECT 1385.395 938.500 1385.910 938.640 ;
        RECT 1385.590 938.440 1385.910 938.500 ;
        RECT 1385.590 917.700 1385.910 917.960 ;
        RECT 1385.680 917.220 1385.820 917.700 ;
        RECT 1386.050 917.220 1386.370 917.280 ;
        RECT 1385.680 917.080 1386.370 917.220 ;
        RECT 1386.050 917.020 1386.370 917.080 ;
        RECT 1386.050 890.020 1386.370 890.080 ;
        RECT 1386.970 890.020 1387.290 890.080 ;
        RECT 1386.050 889.880 1387.290 890.020 ;
        RECT 1386.050 889.820 1386.370 889.880 ;
        RECT 1386.970 889.820 1387.290 889.880 ;
        RECT 1385.590 800.600 1385.910 800.660 ;
        RECT 1386.970 800.600 1387.290 800.660 ;
        RECT 1385.590 800.460 1387.290 800.600 ;
        RECT 1385.590 800.400 1385.910 800.460 ;
        RECT 1386.970 800.400 1387.290 800.460 ;
        RECT 1385.590 793.460 1385.910 793.520 ;
        RECT 1386.050 793.460 1386.370 793.520 ;
        RECT 1385.590 793.320 1386.370 793.460 ;
        RECT 1385.590 793.260 1385.910 793.320 ;
        RECT 1386.050 793.260 1386.370 793.320 ;
        RECT 1385.590 745.180 1385.910 745.240 ;
        RECT 1385.395 745.040 1385.910 745.180 ;
        RECT 1385.590 744.980 1385.910 745.040 ;
        RECT 1385.605 697.240 1385.895 697.285 ;
        RECT 1386.050 697.240 1386.370 697.300 ;
        RECT 1385.605 697.100 1386.370 697.240 ;
        RECT 1385.605 697.055 1385.895 697.100 ;
        RECT 1386.050 697.040 1386.370 697.100 ;
        RECT 1386.050 579.940 1386.370 580.000 ;
        RECT 1385.855 579.800 1386.370 579.940 ;
        RECT 1386.050 579.740 1386.370 579.800 ;
        RECT 1386.050 511.260 1386.370 511.320 ;
        RECT 1385.855 511.120 1386.370 511.260 ;
        RECT 1386.050 511.060 1386.370 511.120 ;
        RECT 1384.670 455.500 1384.990 455.560 ;
        RECT 1385.590 455.500 1385.910 455.560 ;
        RECT 1384.670 455.360 1385.910 455.500 ;
        RECT 1384.670 455.300 1384.990 455.360 ;
        RECT 1385.590 455.300 1385.910 455.360 ;
        RECT 1385.590 420.820 1385.910 420.880 ;
        RECT 1385.395 420.680 1385.910 420.820 ;
        RECT 1385.590 420.620 1385.910 420.680 ;
        RECT 1385.590 372.880 1385.910 372.940 ;
        RECT 1385.395 372.740 1385.910 372.880 ;
        RECT 1385.590 372.680 1385.910 372.740 ;
        RECT 1385.590 365.400 1385.910 365.460 ;
        RECT 1385.395 365.260 1385.910 365.400 ;
        RECT 1385.590 365.200 1385.910 365.260 ;
        RECT 1385.605 317.800 1385.895 317.845 ;
        RECT 1386.050 317.800 1386.370 317.860 ;
        RECT 1385.605 317.660 1386.370 317.800 ;
        RECT 1385.605 317.615 1385.895 317.660 ;
        RECT 1386.050 317.600 1386.370 317.660 ;
        RECT 1385.590 241.640 1385.910 241.700 ;
        RECT 1386.050 241.640 1386.370 241.700 ;
        RECT 1385.590 241.500 1386.370 241.640 ;
        RECT 1385.590 241.440 1385.910 241.500 ;
        RECT 1386.050 241.440 1386.370 241.500 ;
        RECT 1385.590 17.580 1385.910 17.640 ;
        RECT 2286.270 17.580 2286.590 17.640 ;
        RECT 1385.590 17.440 2286.590 17.580 ;
        RECT 1385.590 17.380 1385.910 17.440 ;
        RECT 2286.270 17.380 2286.590 17.440 ;
      LAYER via ;
        RECT 1385.160 1692.560 1385.420 1692.820 ;
        RECT 1385.160 1676.920 1385.420 1677.180 ;
        RECT 1385.160 1635.100 1385.420 1635.360 ;
        RECT 1385.620 1635.100 1385.880 1635.360 ;
        RECT 1385.620 1452.180 1385.880 1452.440 ;
        RECT 1386.540 1452.180 1386.800 1452.440 ;
        RECT 1385.620 1448.780 1385.880 1449.040 ;
        RECT 1386.540 1448.780 1386.800 1449.040 ;
        RECT 1386.080 1372.960 1386.340 1373.220 ;
        RECT 1386.080 1324.680 1386.340 1324.940 ;
        RECT 1386.080 1276.060 1386.340 1276.320 ;
        RECT 1386.080 1234.920 1386.340 1235.180 ;
        RECT 1386.080 1207.380 1386.340 1207.640 ;
        RECT 1386.080 1186.980 1386.340 1187.240 ;
        RECT 1385.620 1048.600 1385.880 1048.860 ;
        RECT 1386.080 1048.600 1386.340 1048.860 ;
        RECT 1385.620 1041.460 1385.880 1041.720 ;
        RECT 1386.080 1041.460 1386.340 1041.720 ;
        RECT 1385.620 986.380 1385.880 986.640 ;
        RECT 1385.620 938.440 1385.880 938.700 ;
        RECT 1385.620 917.700 1385.880 917.960 ;
        RECT 1386.080 917.020 1386.340 917.280 ;
        RECT 1386.080 889.820 1386.340 890.080 ;
        RECT 1387.000 889.820 1387.260 890.080 ;
        RECT 1385.620 800.400 1385.880 800.660 ;
        RECT 1387.000 800.400 1387.260 800.660 ;
        RECT 1385.620 793.260 1385.880 793.520 ;
        RECT 1386.080 793.260 1386.340 793.520 ;
        RECT 1385.620 744.980 1385.880 745.240 ;
        RECT 1386.080 697.040 1386.340 697.300 ;
        RECT 1386.080 579.740 1386.340 580.000 ;
        RECT 1386.080 511.060 1386.340 511.320 ;
        RECT 1384.700 455.300 1384.960 455.560 ;
        RECT 1385.620 455.300 1385.880 455.560 ;
        RECT 1385.620 420.620 1385.880 420.880 ;
        RECT 1385.620 372.680 1385.880 372.940 ;
        RECT 1385.620 365.200 1385.880 365.460 ;
        RECT 1386.080 317.600 1386.340 317.860 ;
        RECT 1385.620 241.440 1385.880 241.700 ;
        RECT 1386.080 241.440 1386.340 241.700 ;
        RECT 1385.620 17.380 1385.880 17.640 ;
        RECT 2286.300 17.380 2286.560 17.640 ;
      LAYER met2 ;
        RECT 1384.600 1700.410 1384.880 1704.000 ;
        RECT 1384.600 1700.270 1385.360 1700.410 ;
        RECT 1384.600 1700.000 1384.880 1700.270 ;
        RECT 1385.220 1692.850 1385.360 1700.270 ;
        RECT 1385.160 1692.530 1385.420 1692.850 ;
        RECT 1385.160 1676.890 1385.420 1677.210 ;
        RECT 1385.220 1635.390 1385.360 1676.890 ;
        RECT 1385.160 1635.070 1385.420 1635.390 ;
        RECT 1385.620 1635.070 1385.880 1635.390 ;
        RECT 1385.680 1563.050 1385.820 1635.070 ;
        RECT 1385.680 1562.910 1386.740 1563.050 ;
        RECT 1386.600 1452.470 1386.740 1562.910 ;
        RECT 1385.620 1452.150 1385.880 1452.470 ;
        RECT 1386.540 1452.150 1386.800 1452.470 ;
        RECT 1385.680 1449.070 1385.820 1452.150 ;
        RECT 1385.620 1448.750 1385.880 1449.070 ;
        RECT 1386.540 1448.750 1386.800 1449.070 ;
        RECT 1386.600 1417.530 1386.740 1448.750 ;
        RECT 1386.140 1417.390 1386.740 1417.530 ;
        RECT 1386.140 1373.250 1386.280 1417.390 ;
        RECT 1386.080 1372.930 1386.340 1373.250 ;
        RECT 1386.080 1324.650 1386.340 1324.970 ;
        RECT 1386.140 1276.350 1386.280 1324.650 ;
        RECT 1386.080 1276.030 1386.340 1276.350 ;
        RECT 1386.080 1234.890 1386.340 1235.210 ;
        RECT 1386.140 1207.670 1386.280 1234.890 ;
        RECT 1386.080 1207.350 1386.340 1207.670 ;
        RECT 1386.080 1186.950 1386.340 1187.270 ;
        RECT 1386.140 1048.890 1386.280 1186.950 ;
        RECT 1385.620 1048.570 1385.880 1048.890 ;
        RECT 1386.080 1048.570 1386.340 1048.890 ;
        RECT 1385.680 1041.750 1385.820 1048.570 ;
        RECT 1385.620 1041.430 1385.880 1041.750 ;
        RECT 1386.080 1041.430 1386.340 1041.750 ;
        RECT 1386.140 993.890 1386.280 1041.430 ;
        RECT 1385.680 993.750 1386.280 993.890 ;
        RECT 1385.680 986.670 1385.820 993.750 ;
        RECT 1385.620 986.350 1385.880 986.670 ;
        RECT 1385.620 938.410 1385.880 938.730 ;
        RECT 1385.680 917.990 1385.820 938.410 ;
        RECT 1385.620 917.670 1385.880 917.990 ;
        RECT 1386.080 916.990 1386.340 917.310 ;
        RECT 1386.140 890.110 1386.280 916.990 ;
        RECT 1386.080 889.790 1386.340 890.110 ;
        RECT 1387.000 889.790 1387.260 890.110 ;
        RECT 1387.060 800.690 1387.200 889.790 ;
        RECT 1385.620 800.370 1385.880 800.690 ;
        RECT 1387.000 800.370 1387.260 800.690 ;
        RECT 1385.680 793.550 1385.820 800.370 ;
        RECT 1385.620 793.230 1385.880 793.550 ;
        RECT 1386.080 793.230 1386.340 793.550 ;
        RECT 1386.140 745.690 1386.280 793.230 ;
        RECT 1385.680 745.550 1386.280 745.690 ;
        RECT 1385.680 745.270 1385.820 745.550 ;
        RECT 1385.620 744.950 1385.880 745.270 ;
        RECT 1386.080 697.010 1386.340 697.330 ;
        RECT 1386.140 580.030 1386.280 697.010 ;
        RECT 1386.080 579.710 1386.340 580.030 ;
        RECT 1386.080 511.030 1386.340 511.350 ;
        RECT 1386.140 503.725 1386.280 511.030 ;
        RECT 1384.690 503.355 1384.970 503.725 ;
        RECT 1386.070 503.355 1386.350 503.725 ;
        RECT 1384.760 455.590 1384.900 503.355 ;
        RECT 1384.700 455.270 1384.960 455.590 ;
        RECT 1385.620 455.270 1385.880 455.590 ;
        RECT 1385.680 420.910 1385.820 455.270 ;
        RECT 1385.620 420.590 1385.880 420.910 ;
        RECT 1385.620 372.650 1385.880 372.970 ;
        RECT 1385.680 365.490 1385.820 372.650 ;
        RECT 1385.620 365.170 1385.880 365.490 ;
        RECT 1386.080 317.570 1386.340 317.890 ;
        RECT 1386.140 241.730 1386.280 317.570 ;
        RECT 1385.620 241.410 1385.880 241.730 ;
        RECT 1386.080 241.410 1386.340 241.730 ;
        RECT 1385.680 17.670 1385.820 241.410 ;
        RECT 1385.620 17.350 1385.880 17.670 ;
        RECT 2286.300 17.350 2286.560 17.670 ;
        RECT 2286.360 2.400 2286.500 17.350 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
      LAYER via2 ;
        RECT 1384.690 503.400 1384.970 503.680 ;
        RECT 1386.070 503.400 1386.350 503.680 ;
      LAYER met3 ;
        RECT 1384.665 503.690 1384.995 503.705 ;
        RECT 1386.045 503.690 1386.375 503.705 ;
        RECT 1384.665 503.390 1386.375 503.690 ;
        RECT 1384.665 503.375 1384.995 503.390 ;
        RECT 1386.045 503.375 1386.375 503.390 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1386.585 1621.545 1386.755 1656.395 ;
        RECT 1385.205 1283.585 1385.375 1331.695 ;
        RECT 1384.745 1248.565 1384.915 1283.415 ;
        RECT 1384.745 510.765 1384.915 558.875 ;
        RECT 1384.285 186.405 1384.455 224.995 ;
      LAYER mcon ;
        RECT 1386.585 1656.225 1386.755 1656.395 ;
        RECT 1385.205 1331.525 1385.375 1331.695 ;
        RECT 1384.745 1283.245 1384.915 1283.415 ;
        RECT 1384.745 558.705 1384.915 558.875 ;
        RECT 1384.285 224.825 1384.455 224.995 ;
      LAYER met1 ;
        RECT 1385.130 1686.300 1385.450 1686.360 ;
        RECT 1386.970 1686.300 1387.290 1686.360 ;
        RECT 1385.130 1686.160 1387.290 1686.300 ;
        RECT 1385.130 1686.100 1385.450 1686.160 ;
        RECT 1386.970 1686.100 1387.290 1686.160 ;
        RECT 1386.510 1656.380 1386.830 1656.440 ;
        RECT 1386.315 1656.240 1386.830 1656.380 ;
        RECT 1386.510 1656.180 1386.830 1656.240 ;
        RECT 1386.525 1621.700 1386.815 1621.745 ;
        RECT 1386.970 1621.700 1387.290 1621.760 ;
        RECT 1386.525 1621.560 1387.290 1621.700 ;
        RECT 1386.525 1621.515 1386.815 1621.560 ;
        RECT 1386.970 1621.500 1387.290 1621.560 ;
        RECT 1385.130 1418.040 1385.450 1418.100 ;
        RECT 1386.050 1418.040 1386.370 1418.100 ;
        RECT 1385.130 1417.900 1386.370 1418.040 ;
        RECT 1385.130 1417.840 1385.450 1417.900 ;
        RECT 1386.050 1417.840 1386.370 1417.900 ;
        RECT 1384.670 1331.680 1384.990 1331.740 ;
        RECT 1385.145 1331.680 1385.435 1331.725 ;
        RECT 1384.670 1331.540 1385.435 1331.680 ;
        RECT 1384.670 1331.480 1384.990 1331.540 ;
        RECT 1385.145 1331.495 1385.435 1331.540 ;
        RECT 1385.130 1283.740 1385.450 1283.800 ;
        RECT 1384.935 1283.600 1385.450 1283.740 ;
        RECT 1385.130 1283.540 1385.450 1283.600 ;
        RECT 1384.670 1283.400 1384.990 1283.460 ;
        RECT 1384.475 1283.260 1384.990 1283.400 ;
        RECT 1384.670 1283.200 1384.990 1283.260 ;
        RECT 1384.670 1248.720 1384.990 1248.780 ;
        RECT 1384.475 1248.580 1384.990 1248.720 ;
        RECT 1384.670 1248.520 1384.990 1248.580 ;
        RECT 1384.670 1145.360 1384.990 1145.420 ;
        RECT 1385.130 1145.360 1385.450 1145.420 ;
        RECT 1384.670 1145.220 1385.450 1145.360 ;
        RECT 1384.670 1145.160 1384.990 1145.220 ;
        RECT 1385.130 1145.160 1385.450 1145.220 ;
        RECT 1384.670 917.900 1384.990 917.960 ;
        RECT 1385.130 917.900 1385.450 917.960 ;
        RECT 1384.670 917.760 1385.450 917.900 ;
        RECT 1384.670 917.700 1384.990 917.760 ;
        RECT 1385.130 917.700 1385.450 917.760 ;
        RECT 1384.210 800.600 1384.530 800.660 ;
        RECT 1385.130 800.600 1385.450 800.660 ;
        RECT 1384.210 800.460 1385.450 800.600 ;
        RECT 1384.210 800.400 1384.530 800.460 ;
        RECT 1385.130 800.400 1385.450 800.460 ;
        RECT 1384.670 662.560 1384.990 662.620 ;
        RECT 1385.130 662.560 1385.450 662.620 ;
        RECT 1384.670 662.420 1385.450 662.560 ;
        RECT 1384.670 662.360 1384.990 662.420 ;
        RECT 1385.130 662.360 1385.450 662.420 ;
        RECT 1384.670 558.860 1384.990 558.920 ;
        RECT 1384.475 558.720 1384.990 558.860 ;
        RECT 1384.670 558.660 1384.990 558.720 ;
        RECT 1384.685 510.920 1384.975 510.965 ;
        RECT 1385.130 510.920 1385.450 510.980 ;
        RECT 1384.685 510.780 1385.450 510.920 ;
        RECT 1384.685 510.735 1384.975 510.780 ;
        RECT 1385.130 510.720 1385.450 510.780 ;
        RECT 1384.670 269.180 1384.990 269.240 ;
        RECT 1385.130 269.180 1385.450 269.240 ;
        RECT 1384.670 269.040 1385.450 269.180 ;
        RECT 1384.670 268.980 1384.990 269.040 ;
        RECT 1385.130 268.980 1385.450 269.040 ;
        RECT 1384.225 224.980 1384.515 225.025 ;
        RECT 1384.670 224.980 1384.990 225.040 ;
        RECT 1384.225 224.840 1384.990 224.980 ;
        RECT 1384.225 224.795 1384.515 224.840 ;
        RECT 1384.670 224.780 1384.990 224.840 ;
        RECT 1384.210 186.560 1384.530 186.620 ;
        RECT 1384.015 186.420 1384.530 186.560 ;
        RECT 1384.210 186.360 1384.530 186.420 ;
        RECT 1384.210 17.240 1384.530 17.300 ;
        RECT 2304.210 17.240 2304.530 17.300 ;
        RECT 1384.210 17.100 2304.530 17.240 ;
        RECT 1384.210 17.040 1384.530 17.100 ;
        RECT 2304.210 17.040 2304.530 17.100 ;
      LAYER via ;
        RECT 1385.160 1686.100 1385.420 1686.360 ;
        RECT 1387.000 1686.100 1387.260 1686.360 ;
        RECT 1386.540 1656.180 1386.800 1656.440 ;
        RECT 1387.000 1621.500 1387.260 1621.760 ;
        RECT 1385.160 1417.840 1385.420 1418.100 ;
        RECT 1386.080 1417.840 1386.340 1418.100 ;
        RECT 1384.700 1331.480 1384.960 1331.740 ;
        RECT 1385.160 1283.540 1385.420 1283.800 ;
        RECT 1384.700 1283.200 1384.960 1283.460 ;
        RECT 1384.700 1248.520 1384.960 1248.780 ;
        RECT 1384.700 1145.160 1384.960 1145.420 ;
        RECT 1385.160 1145.160 1385.420 1145.420 ;
        RECT 1384.700 917.700 1384.960 917.960 ;
        RECT 1385.160 917.700 1385.420 917.960 ;
        RECT 1384.240 800.400 1384.500 800.660 ;
        RECT 1385.160 800.400 1385.420 800.660 ;
        RECT 1384.700 662.360 1384.960 662.620 ;
        RECT 1385.160 662.360 1385.420 662.620 ;
        RECT 1384.700 558.660 1384.960 558.920 ;
        RECT 1385.160 510.720 1385.420 510.980 ;
        RECT 1384.700 268.980 1384.960 269.240 ;
        RECT 1385.160 268.980 1385.420 269.240 ;
        RECT 1384.700 224.780 1384.960 225.040 ;
        RECT 1384.240 186.360 1384.500 186.620 ;
        RECT 1384.240 17.040 1384.500 17.300 ;
        RECT 2304.240 17.040 2304.500 17.300 ;
      LAYER met2 ;
        RECT 1386.440 1700.410 1386.720 1704.000 ;
        RECT 1386.440 1700.270 1387.200 1700.410 ;
        RECT 1386.440 1700.000 1386.720 1700.270 ;
        RECT 1387.060 1686.390 1387.200 1700.270 ;
        RECT 1385.160 1686.070 1385.420 1686.390 ;
        RECT 1387.000 1686.070 1387.260 1686.390 ;
        RECT 1385.220 1678.085 1385.360 1686.070 ;
        RECT 1385.150 1677.715 1385.430 1678.085 ;
        RECT 1386.530 1676.525 1386.810 1676.895 ;
        RECT 1386.600 1656.470 1386.740 1676.525 ;
        RECT 1386.540 1656.150 1386.800 1656.470 ;
        RECT 1387.000 1621.645 1387.260 1621.790 ;
        RECT 1385.150 1621.275 1385.430 1621.645 ;
        RECT 1386.990 1621.275 1387.270 1621.645 ;
        RECT 1385.220 1486.890 1385.360 1621.275 ;
        RECT 1385.220 1486.750 1386.280 1486.890 ;
        RECT 1386.140 1418.130 1386.280 1486.750 ;
        RECT 1385.160 1417.810 1385.420 1418.130 ;
        RECT 1386.080 1417.810 1386.340 1418.130 ;
        RECT 1385.220 1380.245 1385.360 1417.810 ;
        RECT 1384.230 1379.875 1384.510 1380.245 ;
        RECT 1385.150 1379.875 1385.430 1380.245 ;
        RECT 1384.300 1355.650 1384.440 1379.875 ;
        RECT 1384.300 1355.510 1384.900 1355.650 ;
        RECT 1384.760 1331.770 1384.900 1355.510 ;
        RECT 1384.700 1331.450 1384.960 1331.770 ;
        RECT 1385.160 1283.570 1385.420 1283.830 ;
        RECT 1384.760 1283.510 1385.420 1283.570 ;
        RECT 1384.760 1283.490 1385.360 1283.510 ;
        RECT 1384.700 1283.430 1385.360 1283.490 ;
        RECT 1384.700 1283.170 1384.960 1283.430 ;
        RECT 1384.700 1248.490 1384.960 1248.810 ;
        RECT 1384.760 1235.290 1384.900 1248.490 ;
        RECT 1384.760 1235.150 1385.360 1235.290 ;
        RECT 1385.220 1145.450 1385.360 1235.150 ;
        RECT 1384.700 1145.130 1384.960 1145.450 ;
        RECT 1385.160 1145.130 1385.420 1145.450 ;
        RECT 1384.760 1000.010 1384.900 1145.130 ;
        RECT 1384.760 999.870 1385.360 1000.010 ;
        RECT 1385.220 976.210 1385.360 999.870 ;
        RECT 1384.300 976.070 1385.360 976.210 ;
        RECT 1384.300 952.410 1384.440 976.070 ;
        RECT 1384.300 952.270 1384.900 952.410 ;
        RECT 1384.760 917.990 1384.900 952.270 ;
        RECT 1384.700 917.670 1384.960 917.990 ;
        RECT 1385.160 917.670 1385.420 917.990 ;
        RECT 1385.220 879.650 1385.360 917.670 ;
        RECT 1384.760 879.510 1385.360 879.650 ;
        RECT 1384.760 824.570 1384.900 879.510 ;
        RECT 1384.300 824.430 1384.900 824.570 ;
        RECT 1384.300 800.690 1384.440 824.430 ;
        RECT 1384.240 800.370 1384.500 800.690 ;
        RECT 1385.160 800.370 1385.420 800.690 ;
        RECT 1385.220 662.650 1385.360 800.370 ;
        RECT 1384.700 662.330 1384.960 662.650 ;
        RECT 1385.160 662.330 1385.420 662.650 ;
        RECT 1384.760 558.950 1384.900 662.330 ;
        RECT 1384.700 558.630 1384.960 558.950 ;
        RECT 1385.160 510.690 1385.420 511.010 ;
        RECT 1385.220 342.450 1385.360 510.690 ;
        RECT 1384.760 342.310 1385.360 342.450 ;
        RECT 1384.760 341.090 1384.900 342.310 ;
        RECT 1384.760 340.950 1385.360 341.090 ;
        RECT 1385.220 269.270 1385.360 340.950 ;
        RECT 1384.700 268.950 1384.960 269.270 ;
        RECT 1385.160 268.950 1385.420 269.270 ;
        RECT 1384.760 225.070 1384.900 268.950 ;
        RECT 1384.700 224.750 1384.960 225.070 ;
        RECT 1384.240 186.330 1384.500 186.650 ;
        RECT 1384.300 165.650 1384.440 186.330 ;
        RECT 1384.300 165.510 1384.900 165.650 ;
        RECT 1384.760 99.010 1384.900 165.510 ;
        RECT 1383.840 98.870 1384.900 99.010 ;
        RECT 1383.840 96.290 1383.980 98.870 ;
        RECT 1383.840 96.150 1384.440 96.290 ;
        RECT 1384.300 17.330 1384.440 96.150 ;
        RECT 1384.240 17.010 1384.500 17.330 ;
        RECT 2304.240 17.010 2304.500 17.330 ;
        RECT 2304.300 2.400 2304.440 17.010 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
      LAYER via2 ;
        RECT 1385.150 1677.760 1385.430 1678.040 ;
        RECT 1386.530 1676.570 1386.810 1676.850 ;
        RECT 1385.150 1621.320 1385.430 1621.600 ;
        RECT 1386.990 1621.320 1387.270 1621.600 ;
        RECT 1384.230 1379.920 1384.510 1380.200 ;
        RECT 1385.150 1379.920 1385.430 1380.200 ;
      LAYER met3 ;
        RECT 1385.125 1678.050 1385.455 1678.065 ;
        RECT 1385.125 1677.750 1386.130 1678.050 ;
        RECT 1385.125 1677.735 1385.455 1677.750 ;
        RECT 1385.830 1676.860 1386.130 1677.750 ;
        RECT 1386.505 1676.860 1386.835 1676.875 ;
        RECT 1385.830 1676.560 1386.835 1676.860 ;
        RECT 1386.505 1676.545 1386.835 1676.560 ;
        RECT 1385.125 1621.610 1385.455 1621.625 ;
        RECT 1386.965 1621.610 1387.295 1621.625 ;
        RECT 1385.125 1621.310 1387.295 1621.610 ;
        RECT 1385.125 1621.295 1385.455 1621.310 ;
        RECT 1386.965 1621.295 1387.295 1621.310 ;
        RECT 1384.205 1380.210 1384.535 1380.225 ;
        RECT 1385.125 1380.210 1385.455 1380.225 ;
        RECT 1384.205 1379.910 1385.455 1380.210 ;
        RECT 1384.205 1379.895 1384.535 1379.910 ;
        RECT 1385.125 1379.895 1385.455 1379.910 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1388.810 1550.640 1389.130 1550.700 ;
        RECT 1389.730 1550.640 1390.050 1550.700 ;
        RECT 1388.810 1550.500 1390.050 1550.640 ;
        RECT 1388.810 1550.440 1389.130 1550.500 ;
        RECT 1389.730 1550.440 1390.050 1550.500 ;
        RECT 1388.810 1510.860 1389.130 1510.920 ;
        RECT 1389.730 1510.860 1390.050 1510.920 ;
        RECT 1388.810 1510.720 1390.050 1510.860 ;
        RECT 1388.810 1510.660 1389.130 1510.720 ;
        RECT 1389.730 1510.660 1390.050 1510.720 ;
        RECT 1387.890 1063.760 1388.210 1063.820 ;
        RECT 1389.730 1063.760 1390.050 1063.820 ;
        RECT 1387.890 1063.620 1390.050 1063.760 ;
        RECT 1387.890 1063.560 1388.210 1063.620 ;
        RECT 1389.730 1063.560 1390.050 1063.620 ;
        RECT 1388.810 979.580 1389.130 979.840 ;
        RECT 1388.900 979.440 1389.040 979.580 ;
        RECT 1389.730 979.440 1390.050 979.500 ;
        RECT 1388.900 979.300 1390.050 979.440 ;
        RECT 1389.730 979.240 1390.050 979.300 ;
        RECT 1387.890 302.160 1388.210 302.220 ;
        RECT 1389.730 302.160 1390.050 302.220 ;
        RECT 1387.890 302.020 1390.050 302.160 ;
        RECT 1387.890 301.960 1388.210 302.020 ;
        RECT 1389.730 301.960 1390.050 302.020 ;
        RECT 1388.810 206.760 1389.130 207.020 ;
        RECT 1388.900 206.620 1389.040 206.760 ;
        RECT 1389.730 206.620 1390.050 206.680 ;
        RECT 1388.900 206.480 1390.050 206.620 ;
        RECT 1389.730 206.420 1390.050 206.480 ;
        RECT 1388.810 110.740 1389.130 110.800 ;
        RECT 1389.730 110.740 1390.050 110.800 ;
        RECT 1388.810 110.600 1390.050 110.740 ;
        RECT 1388.810 110.540 1389.130 110.600 ;
        RECT 1389.730 110.540 1390.050 110.600 ;
        RECT 1388.810 86.260 1389.130 86.320 ;
        RECT 1390.650 86.260 1390.970 86.320 ;
        RECT 1388.810 86.120 1390.970 86.260 ;
        RECT 1388.810 86.060 1389.130 86.120 ;
        RECT 1390.650 86.060 1390.970 86.120 ;
      LAYER via ;
        RECT 1388.840 1550.440 1389.100 1550.700 ;
        RECT 1389.760 1550.440 1390.020 1550.700 ;
        RECT 1388.840 1510.660 1389.100 1510.920 ;
        RECT 1389.760 1510.660 1390.020 1510.920 ;
        RECT 1387.920 1063.560 1388.180 1063.820 ;
        RECT 1389.760 1063.560 1390.020 1063.820 ;
        RECT 1388.840 979.580 1389.100 979.840 ;
        RECT 1389.760 979.240 1390.020 979.500 ;
        RECT 1387.920 301.960 1388.180 302.220 ;
        RECT 1389.760 301.960 1390.020 302.220 ;
        RECT 1388.840 206.760 1389.100 207.020 ;
        RECT 1389.760 206.420 1390.020 206.680 ;
        RECT 1388.840 110.540 1389.100 110.800 ;
        RECT 1389.760 110.540 1390.020 110.800 ;
        RECT 1388.840 86.060 1389.100 86.320 ;
        RECT 1390.680 86.060 1390.940 86.320 ;
      LAYER met2 ;
        RECT 1388.280 1700.410 1388.560 1704.000 ;
        RECT 1388.280 1700.270 1389.040 1700.410 ;
        RECT 1388.280 1700.000 1388.560 1700.270 ;
        RECT 1388.900 1667.090 1389.040 1700.270 ;
        RECT 1388.900 1666.950 1389.960 1667.090 ;
        RECT 1389.820 1550.730 1389.960 1666.950 ;
        RECT 1388.840 1550.410 1389.100 1550.730 ;
        RECT 1389.760 1550.410 1390.020 1550.730 ;
        RECT 1388.900 1510.950 1389.040 1550.410 ;
        RECT 1388.840 1510.630 1389.100 1510.950 ;
        RECT 1389.760 1510.630 1390.020 1510.950 ;
        RECT 1389.820 1063.850 1389.960 1510.630 ;
        RECT 1387.920 1063.530 1388.180 1063.850 ;
        RECT 1389.760 1063.530 1390.020 1063.850 ;
        RECT 1387.980 1062.685 1388.120 1063.530 ;
        RECT 1387.910 1062.315 1388.190 1062.685 ;
        RECT 1388.830 1062.315 1389.110 1062.685 ;
        RECT 1388.900 979.870 1389.040 1062.315 ;
        RECT 1388.840 979.550 1389.100 979.870 ;
        RECT 1389.760 979.210 1390.020 979.530 ;
        RECT 1389.820 302.250 1389.960 979.210 ;
        RECT 1387.920 301.930 1388.180 302.250 ;
        RECT 1389.760 301.930 1390.020 302.250 ;
        RECT 1387.980 265.610 1388.120 301.930 ;
        RECT 1387.980 265.470 1389.040 265.610 ;
        RECT 1388.900 207.050 1389.040 265.470 ;
        RECT 1388.840 206.730 1389.100 207.050 ;
        RECT 1389.760 206.390 1390.020 206.710 ;
        RECT 1389.820 110.830 1389.960 206.390 ;
        RECT 1388.840 110.510 1389.100 110.830 ;
        RECT 1389.760 110.510 1390.020 110.830 ;
        RECT 1388.900 86.350 1389.040 110.510 ;
        RECT 1388.840 86.030 1389.100 86.350 ;
        RECT 1390.680 86.030 1390.940 86.350 ;
        RECT 1390.740 20.245 1390.880 86.030 ;
        RECT 1390.670 19.875 1390.950 20.245 ;
        RECT 2322.170 19.875 2322.450 20.245 ;
        RECT 2322.240 2.400 2322.380 19.875 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
      LAYER via2 ;
        RECT 1387.910 1062.360 1388.190 1062.640 ;
        RECT 1388.830 1062.360 1389.110 1062.640 ;
        RECT 1390.670 19.920 1390.950 20.200 ;
        RECT 2322.170 19.920 2322.450 20.200 ;
      LAYER met3 ;
        RECT 1387.885 1062.650 1388.215 1062.665 ;
        RECT 1388.805 1062.650 1389.135 1062.665 ;
        RECT 1387.885 1062.350 1389.135 1062.650 ;
        RECT 1387.885 1062.335 1388.215 1062.350 ;
        RECT 1388.805 1062.335 1389.135 1062.350 ;
        RECT 1390.645 20.210 1390.975 20.225 ;
        RECT 2322.145 20.210 2322.475 20.225 ;
        RECT 1390.645 19.910 2322.475 20.210 ;
        RECT 1390.645 19.895 1390.975 19.910 ;
        RECT 2322.145 19.895 2322.475 19.910 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1390.120 1700.340 1390.400 1704.000 ;
        RECT 1390.120 1700.000 1390.420 1700.340 ;
        RECT 1390.280 19.565 1390.420 1700.000 ;
        RECT 1390.210 19.195 1390.490 19.565 ;
        RECT 2339.650 19.195 2339.930 19.565 ;
        RECT 2339.720 2.400 2339.860 19.195 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
      LAYER via2 ;
        RECT 1390.210 19.240 1390.490 19.520 ;
        RECT 2339.650 19.240 2339.930 19.520 ;
      LAYER met3 ;
        RECT 1390.185 19.530 1390.515 19.545 ;
        RECT 2339.625 19.530 2339.955 19.545 ;
        RECT 1390.185 19.230 2339.955 19.530 ;
        RECT 1390.185 19.215 1390.515 19.230 ;
        RECT 2339.625 19.215 2339.955 19.230 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1389.270 1666.580 1389.590 1666.640 ;
        RECT 1392.490 1666.580 1392.810 1666.640 ;
        RECT 1389.270 1666.440 1392.810 1666.580 ;
        RECT 1389.270 1666.380 1389.590 1666.440 ;
        RECT 1392.490 1666.380 1392.810 1666.440 ;
      LAYER via ;
        RECT 1389.300 1666.380 1389.560 1666.640 ;
        RECT 1392.520 1666.380 1392.780 1666.640 ;
      LAYER met2 ;
        RECT 1391.960 1700.340 1392.240 1704.000 ;
        RECT 1391.960 1700.000 1392.260 1700.340 ;
        RECT 1392.120 1684.600 1392.260 1700.000 ;
        RECT 1392.120 1684.460 1392.720 1684.600 ;
        RECT 1392.580 1666.670 1392.720 1684.460 ;
        RECT 1389.300 1666.350 1389.560 1666.670 ;
        RECT 1392.520 1666.350 1392.780 1666.670 ;
        RECT 1389.360 18.885 1389.500 1666.350 ;
        RECT 1389.290 18.515 1389.570 18.885 ;
        RECT 2357.590 18.515 2357.870 18.885 ;
        RECT 2357.660 2.400 2357.800 18.515 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
      LAYER via2 ;
        RECT 1389.290 18.560 1389.570 18.840 ;
        RECT 2357.590 18.560 2357.870 18.840 ;
      LAYER met3 ;
        RECT 1389.265 18.850 1389.595 18.865 ;
        RECT 2357.565 18.850 2357.895 18.865 ;
        RECT 1389.265 18.550 2357.895 18.850 ;
        RECT 1389.265 18.535 1389.595 18.550 ;
        RECT 2357.565 18.535 2357.895 18.550 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1394.790 1630.540 1395.110 1630.600 ;
        RECT 1399.850 1630.540 1400.170 1630.600 ;
        RECT 1394.790 1630.400 1400.170 1630.540 ;
        RECT 1394.790 1630.340 1395.110 1630.400 ;
        RECT 1399.850 1630.340 1400.170 1630.400 ;
        RECT 1399.850 40.160 1400.170 40.420 ;
        RECT 1399.940 39.400 1400.080 40.160 ;
        RECT 1399.850 39.140 1400.170 39.400 ;
      LAYER via ;
        RECT 1394.820 1630.340 1395.080 1630.600 ;
        RECT 1399.880 1630.340 1400.140 1630.600 ;
        RECT 1399.880 40.160 1400.140 40.420 ;
        RECT 1399.880 39.140 1400.140 39.400 ;
      LAYER met2 ;
        RECT 1393.800 1700.410 1394.080 1704.000 ;
        RECT 1393.800 1700.270 1394.560 1700.410 ;
        RECT 1393.800 1700.000 1394.080 1700.270 ;
        RECT 1394.420 1666.410 1394.560 1700.270 ;
        RECT 1394.420 1666.270 1395.020 1666.410 ;
        RECT 1394.880 1630.630 1395.020 1666.270 ;
        RECT 1394.820 1630.310 1395.080 1630.630 ;
        RECT 1399.880 1630.310 1400.140 1630.630 ;
        RECT 1399.940 40.450 1400.080 1630.310 ;
        RECT 1399.880 40.130 1400.140 40.450 ;
        RECT 1399.880 39.110 1400.140 39.430 ;
        RECT 1399.940 18.205 1400.080 39.110 ;
        RECT 1399.870 17.835 1400.150 18.205 ;
        RECT 2375.530 17.835 2375.810 18.205 ;
        RECT 2375.600 2.400 2375.740 17.835 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
      LAYER via2 ;
        RECT 1399.870 17.880 1400.150 18.160 ;
        RECT 2375.530 17.880 2375.810 18.160 ;
      LAYER met3 ;
        RECT 1399.845 18.170 1400.175 18.185 ;
        RECT 2375.505 18.170 2375.835 18.185 ;
        RECT 1399.845 17.870 2375.835 18.170 ;
        RECT 1399.845 17.855 1400.175 17.870 ;
        RECT 2375.505 17.855 2375.835 17.870 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1395.710 1684.260 1396.030 1684.320 ;
        RECT 1400.310 1684.260 1400.630 1684.320 ;
        RECT 1395.710 1684.120 1400.630 1684.260 ;
        RECT 1395.710 1684.060 1396.030 1684.120 ;
        RECT 1400.310 1684.060 1400.630 1684.120 ;
        RECT 1399.390 34.580 1399.710 34.640 ;
        RECT 1400.310 34.580 1400.630 34.640 ;
        RECT 1399.390 34.440 1400.630 34.580 ;
        RECT 1399.390 34.380 1399.710 34.440 ;
        RECT 1400.310 34.380 1400.630 34.440 ;
      LAYER via ;
        RECT 1395.740 1684.060 1396.000 1684.320 ;
        RECT 1400.340 1684.060 1400.600 1684.320 ;
        RECT 1399.420 34.380 1399.680 34.640 ;
        RECT 1400.340 34.380 1400.600 34.640 ;
      LAYER met2 ;
        RECT 1395.640 1700.340 1395.920 1704.000 ;
        RECT 1395.640 1700.000 1395.940 1700.340 ;
        RECT 1395.800 1684.350 1395.940 1700.000 ;
        RECT 1395.740 1684.030 1396.000 1684.350 ;
        RECT 1400.340 1684.030 1400.600 1684.350 ;
        RECT 1400.400 34.670 1400.540 1684.030 ;
        RECT 1399.420 34.350 1399.680 34.670 ;
        RECT 1400.340 34.350 1400.600 34.670 ;
        RECT 1399.480 17.525 1399.620 34.350 ;
        RECT 1399.410 17.155 1399.690 17.525 ;
        RECT 2393.470 17.155 2393.750 17.525 ;
        RECT 2393.540 2.400 2393.680 17.155 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
      LAYER via2 ;
        RECT 1399.410 17.200 1399.690 17.480 ;
        RECT 2393.470 17.200 2393.750 17.480 ;
      LAYER met3 ;
        RECT 1399.385 17.490 1399.715 17.505 ;
        RECT 2393.445 17.490 2393.775 17.505 ;
        RECT 1399.385 17.190 2393.775 17.490 ;
        RECT 1399.385 17.175 1399.715 17.190 ;
        RECT 2393.445 17.175 2393.775 17.190 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1397.550 1683.920 1397.870 1683.980 ;
        RECT 1399.850 1683.920 1400.170 1683.980 ;
        RECT 1397.550 1683.780 1400.170 1683.920 ;
        RECT 1397.550 1683.720 1397.870 1683.780 ;
        RECT 1399.850 1683.720 1400.170 1683.780 ;
      LAYER via ;
        RECT 1397.580 1683.720 1397.840 1683.980 ;
        RECT 1399.880 1683.720 1400.140 1683.980 ;
      LAYER met2 ;
        RECT 1397.480 1700.340 1397.760 1704.000 ;
        RECT 1397.480 1700.000 1397.780 1700.340 ;
        RECT 1397.640 1684.010 1397.780 1700.000 ;
        RECT 1397.580 1683.690 1397.840 1684.010 ;
        RECT 1399.880 1683.690 1400.140 1684.010 ;
        RECT 1399.940 1631.050 1400.080 1683.690 ;
        RECT 1399.480 1630.910 1400.080 1631.050 ;
        RECT 1399.480 1582.770 1399.620 1630.910 ;
        RECT 1399.020 1582.630 1399.620 1582.770 ;
        RECT 1399.020 1535.850 1399.160 1582.630 ;
        RECT 1399.020 1535.710 1399.620 1535.850 ;
        RECT 1399.480 40.530 1399.620 1535.710 ;
        RECT 1399.020 40.390 1399.620 40.530 ;
        RECT 1399.020 16.845 1399.160 40.390 ;
        RECT 1398.950 16.475 1399.230 16.845 ;
        RECT 2411.410 16.475 2411.690 16.845 ;
        RECT 2411.480 2.400 2411.620 16.475 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
      LAYER via2 ;
        RECT 1398.950 16.520 1399.230 16.800 ;
        RECT 2411.410 16.520 2411.690 16.800 ;
      LAYER met3 ;
        RECT 1398.925 16.810 1399.255 16.825 ;
        RECT 2411.385 16.810 2411.715 16.825 ;
        RECT 1398.925 16.510 2411.715 16.810 ;
        RECT 1398.925 16.495 1399.255 16.510 ;
        RECT 2411.385 16.495 2411.715 16.510 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 806.910 1556.080 807.230 1556.140 ;
        RECT 1232.410 1556.080 1232.730 1556.140 ;
        RECT 806.910 1555.940 1232.730 1556.080 ;
        RECT 806.910 1555.880 807.230 1555.940 ;
        RECT 1232.410 1555.880 1232.730 1555.940 ;
      LAYER via ;
        RECT 806.940 1555.880 807.200 1556.140 ;
        RECT 1232.440 1555.880 1232.700 1556.140 ;
      LAYER met2 ;
        RECT 1232.340 1700.340 1232.620 1704.000 ;
        RECT 1232.340 1700.000 1232.640 1700.340 ;
        RECT 1232.500 1556.170 1232.640 1700.000 ;
        RECT 806.940 1555.850 807.200 1556.170 ;
        RECT 1232.440 1555.850 1232.700 1556.170 ;
        RECT 807.000 18.090 807.140 1555.850 ;
        RECT 805.620 17.950 807.140 18.090 ;
        RECT 805.620 2.400 805.760 17.950 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1121.165 23.885 1121.335 25.075 ;
      LAYER mcon ;
        RECT 1121.165 24.905 1121.335 25.075 ;
      LAYER met1 ;
        RECT 1121.105 25.060 1121.395 25.105 ;
        RECT 1146.390 25.060 1146.710 25.120 ;
        RECT 1121.105 24.920 1146.710 25.060 ;
        RECT 1121.105 24.875 1121.395 24.920 ;
        RECT 1146.390 24.860 1146.710 24.920 ;
        RECT 2.830 24.040 3.150 24.100 ;
        RECT 1121.105 24.040 1121.395 24.085 ;
        RECT 2.830 23.900 1121.395 24.040 ;
        RECT 2.830 23.840 3.150 23.900 ;
        RECT 1121.105 23.855 1121.395 23.900 ;
      LAYER via ;
        RECT 1146.420 24.860 1146.680 25.120 ;
        RECT 2.860 23.840 3.120 24.100 ;
      LAYER met2 ;
        RECT 1150.000 1700.410 1150.280 1704.000 ;
        RECT 1146.480 1700.270 1150.280 1700.410 ;
        RECT 1146.480 25.150 1146.620 1700.270 ;
        RECT 1150.000 1700.000 1150.280 1700.270 ;
        RECT 1146.420 24.830 1146.680 25.150 ;
        RECT 2.860 23.810 3.120 24.130 ;
        RECT 2.920 2.400 3.060 23.810 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 24.380 8.670 24.440 ;
        RECT 8.350 24.240 1121.780 24.380 ;
        RECT 8.350 24.180 8.670 24.240 ;
        RECT 1121.640 24.040 1121.780 24.240 ;
        RECT 1146.850 24.040 1147.170 24.100 ;
        RECT 1121.640 23.900 1147.170 24.040 ;
        RECT 1146.850 23.840 1147.170 23.900 ;
      LAYER via ;
        RECT 8.380 24.180 8.640 24.440 ;
        RECT 1146.880 23.840 1147.140 24.100 ;
      LAYER met2 ;
        RECT 1150.460 1700.340 1150.740 1704.000 ;
        RECT 1150.460 1700.000 1150.760 1700.340 ;
        RECT 1150.620 1677.970 1150.760 1700.000 ;
        RECT 1146.940 1677.830 1150.760 1677.970 ;
        RECT 8.380 24.150 8.640 24.470 ;
        RECT 8.440 2.400 8.580 24.150 ;
        RECT 1146.940 24.130 1147.080 1677.830 ;
        RECT 1146.880 23.810 1147.140 24.130 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1145.930 1678.140 1146.250 1678.200 ;
        RECT 1150.990 1678.140 1151.310 1678.200 ;
        RECT 1145.930 1678.000 1151.310 1678.140 ;
        RECT 1145.930 1677.940 1146.250 1678.000 ;
        RECT 1150.990 1677.940 1151.310 1678.000 ;
        RECT 14.330 24.720 14.650 24.780 ;
        RECT 1145.930 24.720 1146.250 24.780 ;
        RECT 14.330 24.580 1146.250 24.720 ;
        RECT 14.330 24.520 14.650 24.580 ;
        RECT 1145.930 24.520 1146.250 24.580 ;
      LAYER via ;
        RECT 1145.960 1677.940 1146.220 1678.200 ;
        RECT 1151.020 1677.940 1151.280 1678.200 ;
        RECT 14.360 24.520 14.620 24.780 ;
        RECT 1145.960 24.520 1146.220 24.780 ;
      LAYER met2 ;
        RECT 1150.920 1700.340 1151.200 1704.000 ;
        RECT 1150.920 1700.000 1151.220 1700.340 ;
        RECT 1151.080 1678.230 1151.220 1700.000 ;
        RECT 1145.960 1677.910 1146.220 1678.230 ;
        RECT 1151.020 1677.910 1151.280 1678.230 ;
        RECT 1146.020 24.810 1146.160 1677.910 ;
        RECT 14.360 24.490 14.620 24.810 ;
        RECT 1145.960 24.490 1146.220 24.810 ;
        RECT 14.420 2.400 14.560 24.490 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1120.705 22.865 1120.875 25.075 ;
      LAYER mcon ;
        RECT 1120.705 24.905 1120.875 25.075 ;
      LAYER met1 ;
        RECT 38.250 25.060 38.570 25.120 ;
        RECT 1120.645 25.060 1120.935 25.105 ;
        RECT 38.250 24.920 1120.935 25.060 ;
        RECT 38.250 24.860 38.570 24.920 ;
        RECT 1120.645 24.875 1120.935 24.920 ;
        RECT 1120.645 23.020 1120.935 23.065 ;
        RECT 1153.750 23.020 1154.070 23.080 ;
        RECT 1120.645 22.880 1154.070 23.020 ;
        RECT 1120.645 22.835 1120.935 22.880 ;
        RECT 1153.750 22.820 1154.070 22.880 ;
      LAYER via ;
        RECT 38.280 24.860 38.540 25.120 ;
        RECT 1153.780 22.820 1154.040 23.080 ;
      LAYER met2 ;
        RECT 1153.220 1700.410 1153.500 1704.000 ;
        RECT 1153.220 1700.270 1153.980 1700.410 ;
        RECT 1153.220 1700.000 1153.500 1700.270 ;
        RECT 38.280 24.830 38.540 25.150 ;
        RECT 38.340 2.400 38.480 24.830 ;
        RECT 1153.840 23.110 1153.980 1700.270 ;
        RECT 1153.780 22.790 1154.040 23.110 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1168.010 1688.000 1168.330 1688.060 ;
        RECT 1174.450 1688.000 1174.770 1688.060 ;
        RECT 1168.010 1687.860 1174.770 1688.000 ;
        RECT 1168.010 1687.800 1168.330 1687.860 ;
        RECT 1174.450 1687.800 1174.770 1687.860 ;
        RECT 241.110 1680.180 241.430 1680.240 ;
        RECT 1168.010 1680.180 1168.330 1680.240 ;
        RECT 241.110 1680.040 1168.330 1680.180 ;
        RECT 241.110 1679.980 241.430 1680.040 ;
        RECT 1168.010 1679.980 1168.330 1680.040 ;
      LAYER via ;
        RECT 1168.040 1687.800 1168.300 1688.060 ;
        RECT 1174.480 1687.800 1174.740 1688.060 ;
        RECT 241.140 1679.980 241.400 1680.240 ;
        RECT 1168.040 1679.980 1168.300 1680.240 ;
      LAYER met2 ;
        RECT 1174.380 1700.340 1174.660 1704.000 ;
        RECT 1174.380 1700.000 1174.680 1700.340 ;
        RECT 1174.540 1688.090 1174.680 1700.000 ;
        RECT 1168.040 1687.770 1168.300 1688.090 ;
        RECT 1174.480 1687.770 1174.740 1688.090 ;
        RECT 1168.100 1680.270 1168.240 1687.770 ;
        RECT 241.140 1679.950 241.400 1680.270 ;
        RECT 1168.040 1679.950 1168.300 1680.270 ;
        RECT 241.200 17.410 241.340 1679.950 ;
        RECT 240.740 17.270 241.340 17.410 ;
        RECT 240.740 2.400 240.880 17.270 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1159.270 1687.320 1159.590 1687.380 ;
        RECT 1176.290 1687.320 1176.610 1687.380 ;
        RECT 1159.270 1687.180 1176.610 1687.320 ;
        RECT 1159.270 1687.120 1159.590 1687.180 ;
        RECT 1176.290 1687.120 1176.610 1687.180 ;
        RECT 261.810 1673.040 262.130 1673.100 ;
        RECT 1159.270 1673.040 1159.590 1673.100 ;
        RECT 261.810 1672.900 1159.590 1673.040 ;
        RECT 261.810 1672.840 262.130 1672.900 ;
        RECT 1159.270 1672.840 1159.590 1672.900 ;
        RECT 258.130 17.920 258.450 17.980 ;
        RECT 261.810 17.920 262.130 17.980 ;
        RECT 258.130 17.780 262.130 17.920 ;
        RECT 258.130 17.720 258.450 17.780 ;
        RECT 261.810 17.720 262.130 17.780 ;
      LAYER via ;
        RECT 1159.300 1687.120 1159.560 1687.380 ;
        RECT 1176.320 1687.120 1176.580 1687.380 ;
        RECT 261.840 1672.840 262.100 1673.100 ;
        RECT 1159.300 1672.840 1159.560 1673.100 ;
        RECT 258.160 17.720 258.420 17.980 ;
        RECT 261.840 17.720 262.100 17.980 ;
      LAYER met2 ;
        RECT 1176.220 1700.340 1176.500 1704.000 ;
        RECT 1176.220 1700.000 1176.520 1700.340 ;
        RECT 1176.380 1687.410 1176.520 1700.000 ;
        RECT 1159.300 1687.090 1159.560 1687.410 ;
        RECT 1176.320 1687.090 1176.580 1687.410 ;
        RECT 1159.360 1673.130 1159.500 1687.090 ;
        RECT 261.840 1672.810 262.100 1673.130 ;
        RECT 1159.300 1672.810 1159.560 1673.130 ;
        RECT 261.900 18.010 262.040 1672.810 ;
        RECT 258.160 17.690 258.420 18.010 ;
        RECT 261.840 17.690 262.100 18.010 ;
        RECT 258.220 2.400 258.360 17.690 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.510 1666.240 282.830 1666.300 ;
        RECT 1178.130 1666.240 1178.450 1666.300 ;
        RECT 282.510 1666.100 1178.450 1666.240 ;
        RECT 282.510 1666.040 282.830 1666.100 ;
        RECT 1178.130 1666.040 1178.450 1666.100 ;
        RECT 276.070 16.900 276.390 16.960 ;
        RECT 282.510 16.900 282.830 16.960 ;
        RECT 276.070 16.760 282.830 16.900 ;
        RECT 276.070 16.700 276.390 16.760 ;
        RECT 282.510 16.700 282.830 16.760 ;
      LAYER via ;
        RECT 282.540 1666.040 282.800 1666.300 ;
        RECT 1178.160 1666.040 1178.420 1666.300 ;
        RECT 276.100 16.700 276.360 16.960 ;
        RECT 282.540 16.700 282.800 16.960 ;
      LAYER met2 ;
        RECT 1178.060 1700.340 1178.340 1704.000 ;
        RECT 1178.060 1700.000 1178.360 1700.340 ;
        RECT 1178.220 1666.330 1178.360 1700.000 ;
        RECT 282.540 1666.010 282.800 1666.330 ;
        RECT 1178.160 1666.010 1178.420 1666.330 ;
        RECT 282.600 16.990 282.740 1666.010 ;
        RECT 276.100 16.670 276.360 16.990 ;
        RECT 282.540 16.670 282.800 16.990 ;
        RECT 276.160 2.400 276.300 16.670 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1179.970 1675.760 1180.290 1675.820 ;
        RECT 1181.810 1675.760 1182.130 1675.820 ;
        RECT 1179.970 1675.620 1182.130 1675.760 ;
        RECT 1179.970 1675.560 1180.290 1675.620 ;
        RECT 1181.810 1675.560 1182.130 1675.620 ;
        RECT 294.010 45.120 294.330 45.180 ;
        RECT 1181.810 45.120 1182.130 45.180 ;
        RECT 294.010 44.980 1182.130 45.120 ;
        RECT 294.010 44.920 294.330 44.980 ;
        RECT 1181.810 44.920 1182.130 44.980 ;
      LAYER via ;
        RECT 1180.000 1675.560 1180.260 1675.820 ;
        RECT 1181.840 1675.560 1182.100 1675.820 ;
        RECT 294.040 44.920 294.300 45.180 ;
        RECT 1181.840 44.920 1182.100 45.180 ;
      LAYER met2 ;
        RECT 1179.900 1700.340 1180.180 1704.000 ;
        RECT 1179.900 1700.000 1180.200 1700.340 ;
        RECT 1180.060 1675.850 1180.200 1700.000 ;
        RECT 1180.000 1675.530 1180.260 1675.850 ;
        RECT 1181.840 1675.530 1182.100 1675.850 ;
        RECT 1181.900 45.210 1182.040 1675.530 ;
        RECT 294.040 44.890 294.300 45.210 ;
        RECT 1181.840 44.890 1182.100 45.210 ;
        RECT 294.100 2.400 294.240 44.890 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1181.810 1678.480 1182.130 1678.540 ;
        RECT 1181.810 1678.340 1182.960 1678.480 ;
        RECT 1181.810 1678.280 1182.130 1678.340 ;
        RECT 1182.820 1678.200 1182.960 1678.340 ;
        RECT 1182.730 1677.940 1183.050 1678.200 ;
        RECT 311.950 45.460 312.270 45.520 ;
        RECT 1182.730 45.460 1183.050 45.520 ;
        RECT 311.950 45.320 1183.050 45.460 ;
        RECT 311.950 45.260 312.270 45.320 ;
        RECT 1182.730 45.260 1183.050 45.320 ;
      LAYER via ;
        RECT 1181.840 1678.280 1182.100 1678.540 ;
        RECT 1182.760 1677.940 1183.020 1678.200 ;
        RECT 311.980 45.260 312.240 45.520 ;
        RECT 1182.760 45.260 1183.020 45.520 ;
      LAYER met2 ;
        RECT 1181.740 1700.340 1182.020 1704.000 ;
        RECT 1181.740 1700.000 1182.040 1700.340 ;
        RECT 1181.900 1678.570 1182.040 1700.000 ;
        RECT 1181.840 1678.250 1182.100 1678.570 ;
        RECT 1182.760 1677.910 1183.020 1678.230 ;
        RECT 1182.820 45.550 1182.960 1677.910 ;
        RECT 311.980 45.230 312.240 45.550 ;
        RECT 1182.760 45.230 1183.020 45.550 ;
        RECT 312.040 2.400 312.180 45.230 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1182.270 1679.160 1182.590 1679.220 ;
        RECT 1183.190 1679.160 1183.510 1679.220 ;
        RECT 1182.270 1679.020 1183.510 1679.160 ;
        RECT 1182.270 1678.960 1182.590 1679.020 ;
        RECT 1183.190 1678.960 1183.510 1679.020 ;
        RECT 329.890 45.800 330.210 45.860 ;
        RECT 1182.270 45.800 1182.590 45.860 ;
        RECT 329.890 45.660 1182.590 45.800 ;
        RECT 329.890 45.600 330.210 45.660 ;
        RECT 1182.270 45.600 1182.590 45.660 ;
      LAYER via ;
        RECT 1182.300 1678.960 1182.560 1679.220 ;
        RECT 1183.220 1678.960 1183.480 1679.220 ;
        RECT 329.920 45.600 330.180 45.860 ;
        RECT 1182.300 45.600 1182.560 45.860 ;
      LAYER met2 ;
        RECT 1183.580 1700.410 1183.860 1704.000 ;
        RECT 1183.280 1700.270 1183.860 1700.410 ;
        RECT 1183.280 1679.250 1183.420 1700.270 ;
        RECT 1183.580 1700.000 1183.860 1700.270 ;
        RECT 1182.300 1678.930 1182.560 1679.250 ;
        RECT 1183.220 1678.930 1183.480 1679.250 ;
        RECT 1182.360 45.890 1182.500 1678.930 ;
        RECT 329.920 45.570 330.180 45.890 ;
        RECT 1182.300 45.570 1182.560 45.890 ;
        RECT 329.980 2.400 330.120 45.570 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1183.190 1678.140 1183.510 1678.200 ;
        RECT 1185.030 1678.140 1185.350 1678.200 ;
        RECT 1183.190 1678.000 1185.350 1678.140 ;
        RECT 1183.190 1677.940 1183.510 1678.000 ;
        RECT 1185.030 1677.940 1185.350 1678.000 ;
        RECT 347.370 46.140 347.690 46.200 ;
        RECT 1183.190 46.140 1183.510 46.200 ;
        RECT 347.370 46.000 1183.510 46.140 ;
        RECT 347.370 45.940 347.690 46.000 ;
        RECT 1183.190 45.940 1183.510 46.000 ;
      LAYER via ;
        RECT 1183.220 1677.940 1183.480 1678.200 ;
        RECT 1185.060 1677.940 1185.320 1678.200 ;
        RECT 347.400 45.940 347.660 46.200 ;
        RECT 1183.220 45.940 1183.480 46.200 ;
      LAYER met2 ;
        RECT 1185.420 1700.410 1185.700 1704.000 ;
        RECT 1185.120 1700.270 1185.700 1700.410 ;
        RECT 1185.120 1678.230 1185.260 1700.270 ;
        RECT 1185.420 1700.000 1185.700 1700.270 ;
        RECT 1183.220 1677.910 1183.480 1678.230 ;
        RECT 1185.060 1677.910 1185.320 1678.230 ;
        RECT 1183.280 46.230 1183.420 1677.910 ;
        RECT 347.400 45.910 347.660 46.230 ;
        RECT 1183.220 45.910 1183.480 46.230 ;
        RECT 347.460 2.400 347.600 45.910 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 46.480 365.630 46.540 ;
        RECT 1188.250 46.480 1188.570 46.540 ;
        RECT 365.310 46.340 1188.570 46.480 ;
        RECT 365.310 46.280 365.630 46.340 ;
        RECT 1188.250 46.280 1188.570 46.340 ;
      LAYER via ;
        RECT 365.340 46.280 365.600 46.540 ;
        RECT 1188.280 46.280 1188.540 46.540 ;
      LAYER met2 ;
        RECT 1187.260 1700.340 1187.540 1704.000 ;
        RECT 1187.260 1700.000 1187.560 1700.340 ;
        RECT 1187.420 1672.530 1187.560 1700.000 ;
        RECT 1187.420 1672.390 1188.480 1672.530 ;
        RECT 1188.340 46.570 1188.480 1672.390 ;
        RECT 365.340 46.250 365.600 46.570 ;
        RECT 1188.280 46.250 1188.540 46.570 ;
        RECT 365.400 2.400 365.540 46.250 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 46.820 383.570 46.880 ;
        RECT 1188.710 46.820 1189.030 46.880 ;
        RECT 383.250 46.680 1189.030 46.820 ;
        RECT 383.250 46.620 383.570 46.680 ;
        RECT 1188.710 46.620 1189.030 46.680 ;
      LAYER via ;
        RECT 383.280 46.620 383.540 46.880 ;
        RECT 1188.740 46.620 1189.000 46.880 ;
      LAYER met2 ;
        RECT 1189.100 1700.410 1189.380 1704.000 ;
        RECT 1188.800 1700.270 1189.380 1700.410 ;
        RECT 1188.800 46.910 1188.940 1700.270 ;
        RECT 1189.100 1700.000 1189.380 1700.270 ;
        RECT 383.280 46.590 383.540 46.910 ;
        RECT 1188.740 46.590 1189.000 46.910 ;
        RECT 383.340 2.400 383.480 46.590 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 47.160 401.510 47.220 ;
        RECT 1191.010 47.160 1191.330 47.220 ;
        RECT 401.190 47.020 1191.330 47.160 ;
        RECT 401.190 46.960 401.510 47.020 ;
        RECT 1191.010 46.960 1191.330 47.020 ;
      LAYER via ;
        RECT 401.220 46.960 401.480 47.220 ;
        RECT 1191.040 46.960 1191.300 47.220 ;
      LAYER met2 ;
        RECT 1190.940 1700.340 1191.220 1704.000 ;
        RECT 1190.940 1700.000 1191.240 1700.340 ;
        RECT 1191.100 47.250 1191.240 1700.000 ;
        RECT 401.220 46.930 401.480 47.250 ;
        RECT 1191.040 46.930 1191.300 47.250 ;
        RECT 401.280 2.400 401.420 46.930 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1153.290 1678.140 1153.610 1678.200 ;
        RECT 1155.590 1678.140 1155.910 1678.200 ;
        RECT 1153.290 1678.000 1155.910 1678.140 ;
        RECT 1153.290 1677.940 1153.610 1678.000 ;
        RECT 1155.590 1677.940 1155.910 1678.000 ;
        RECT 62.170 30.840 62.490 30.900 ;
        RECT 1153.290 30.840 1153.610 30.900 ;
        RECT 62.170 30.700 1153.610 30.840 ;
        RECT 62.170 30.640 62.490 30.700 ;
        RECT 1153.290 30.640 1153.610 30.700 ;
      LAYER via ;
        RECT 1153.320 1677.940 1153.580 1678.200 ;
        RECT 1155.620 1677.940 1155.880 1678.200 ;
        RECT 62.200 30.640 62.460 30.900 ;
        RECT 1153.320 30.640 1153.580 30.900 ;
      LAYER met2 ;
        RECT 1155.980 1700.410 1156.260 1704.000 ;
        RECT 1155.680 1700.270 1156.260 1700.410 ;
        RECT 1155.680 1678.230 1155.820 1700.270 ;
        RECT 1155.980 1700.000 1156.260 1700.270 ;
        RECT 1153.320 1677.910 1153.580 1678.230 ;
        RECT 1155.620 1677.910 1155.880 1678.230 ;
        RECT 1153.380 30.930 1153.520 1677.910 ;
        RECT 62.200 30.610 62.460 30.930 ;
        RECT 1153.320 30.610 1153.580 30.930 ;
        RECT 62.260 2.400 62.400 30.610 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 47.500 419.450 47.560 ;
        RECT 1192.850 47.500 1193.170 47.560 ;
        RECT 419.130 47.360 1193.170 47.500 ;
        RECT 419.130 47.300 419.450 47.360 ;
        RECT 1192.850 47.300 1193.170 47.360 ;
      LAYER via ;
        RECT 419.160 47.300 419.420 47.560 ;
        RECT 1192.880 47.300 1193.140 47.560 ;
      LAYER met2 ;
        RECT 1192.780 1700.340 1193.060 1704.000 ;
        RECT 1192.780 1700.000 1193.080 1700.340 ;
        RECT 1192.940 47.590 1193.080 1700.000 ;
        RECT 419.160 47.270 419.420 47.590 ;
        RECT 1192.880 47.270 1193.140 47.590 ;
        RECT 419.220 2.400 419.360 47.270 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 436.610 47.840 436.930 47.900 ;
        RECT 1195.150 47.840 1195.470 47.900 ;
        RECT 436.610 47.700 1195.470 47.840 ;
        RECT 436.610 47.640 436.930 47.700 ;
        RECT 1195.150 47.640 1195.470 47.700 ;
      LAYER via ;
        RECT 436.640 47.640 436.900 47.900 ;
        RECT 1195.180 47.640 1195.440 47.900 ;
      LAYER met2 ;
        RECT 1194.620 1700.340 1194.900 1704.000 ;
        RECT 1194.620 1700.000 1194.920 1700.340 ;
        RECT 1194.780 1678.480 1194.920 1700.000 ;
        RECT 1194.780 1678.340 1195.380 1678.480 ;
        RECT 1195.240 47.930 1195.380 1678.340 ;
        RECT 436.640 47.610 436.900 47.930 ;
        RECT 1195.180 47.610 1195.440 47.930 ;
        RECT 436.700 2.400 436.840 47.610 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 454.550 48.180 454.870 48.240 ;
        RECT 1196.070 48.180 1196.390 48.240 ;
        RECT 454.550 48.040 1196.390 48.180 ;
        RECT 454.550 47.980 454.870 48.040 ;
        RECT 1196.070 47.980 1196.390 48.040 ;
      LAYER via ;
        RECT 454.580 47.980 454.840 48.240 ;
        RECT 1196.100 47.980 1196.360 48.240 ;
      LAYER met2 ;
        RECT 1196.460 1700.410 1196.740 1704.000 ;
        RECT 1196.160 1700.270 1196.740 1700.410 ;
        RECT 1196.160 48.270 1196.300 1700.270 ;
        RECT 1196.460 1700.000 1196.740 1700.270 ;
        RECT 454.580 47.950 454.840 48.270 ;
        RECT 1196.100 47.950 1196.360 48.270 ;
        RECT 454.640 2.400 454.780 47.950 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 472.490 44.440 472.810 44.500 ;
        RECT 1198.370 44.440 1198.690 44.500 ;
        RECT 472.490 44.300 1198.690 44.440 ;
        RECT 472.490 44.240 472.810 44.300 ;
        RECT 1198.370 44.240 1198.690 44.300 ;
      LAYER via ;
        RECT 472.520 44.240 472.780 44.500 ;
        RECT 1198.400 44.240 1198.660 44.500 ;
      LAYER met2 ;
        RECT 1198.300 1700.340 1198.580 1704.000 ;
        RECT 1198.300 1700.000 1198.600 1700.340 ;
        RECT 1198.460 44.530 1198.600 1700.000 ;
        RECT 472.520 44.210 472.780 44.530 ;
        RECT 1198.400 44.210 1198.660 44.530 ;
        RECT 472.580 2.400 472.720 44.210 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1195.610 1677.800 1195.930 1677.860 ;
        RECT 1200.210 1677.800 1200.530 1677.860 ;
        RECT 1195.610 1677.660 1200.530 1677.800 ;
        RECT 1195.610 1677.600 1195.930 1677.660 ;
        RECT 1200.210 1677.600 1200.530 1677.660 ;
        RECT 490.430 44.100 490.750 44.160 ;
        RECT 1195.610 44.100 1195.930 44.160 ;
        RECT 490.430 43.960 1195.930 44.100 ;
        RECT 490.430 43.900 490.750 43.960 ;
        RECT 1195.610 43.900 1195.930 43.960 ;
      LAYER via ;
        RECT 1195.640 1677.600 1195.900 1677.860 ;
        RECT 1200.240 1677.600 1200.500 1677.860 ;
        RECT 490.460 43.900 490.720 44.160 ;
        RECT 1195.640 43.900 1195.900 44.160 ;
      LAYER met2 ;
        RECT 1200.140 1700.340 1200.420 1704.000 ;
        RECT 1200.140 1700.000 1200.440 1700.340 ;
        RECT 1200.300 1677.890 1200.440 1700.000 ;
        RECT 1195.640 1677.570 1195.900 1677.890 ;
        RECT 1200.240 1677.570 1200.500 1677.890 ;
        RECT 1195.700 44.190 1195.840 1677.570 ;
        RECT 490.460 43.870 490.720 44.190 ;
        RECT 1195.640 43.870 1195.900 44.190 ;
        RECT 490.520 2.400 490.660 43.870 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.910 43.760 508.230 43.820 ;
        RECT 1202.050 43.760 1202.370 43.820 ;
        RECT 507.910 43.620 1202.370 43.760 ;
        RECT 507.910 43.560 508.230 43.620 ;
        RECT 1202.050 43.560 1202.370 43.620 ;
      LAYER via ;
        RECT 507.940 43.560 508.200 43.820 ;
        RECT 1202.080 43.560 1202.340 43.820 ;
      LAYER met2 ;
        RECT 1201.980 1700.340 1202.260 1704.000 ;
        RECT 1201.980 1700.000 1202.280 1700.340 ;
        RECT 1202.140 43.850 1202.280 1700.000 ;
        RECT 507.940 43.530 508.200 43.850 ;
        RECT 1202.080 43.530 1202.340 43.850 ;
        RECT 508.000 2.400 508.140 43.530 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1201.590 1678.480 1201.910 1678.540 ;
        RECT 1203.890 1678.480 1204.210 1678.540 ;
        RECT 1201.590 1678.340 1204.210 1678.480 ;
        RECT 1201.590 1678.280 1201.910 1678.340 ;
        RECT 1203.890 1678.280 1204.210 1678.340 ;
        RECT 525.850 43.420 526.170 43.480 ;
        RECT 1201.590 43.420 1201.910 43.480 ;
        RECT 525.850 43.280 1201.910 43.420 ;
        RECT 525.850 43.220 526.170 43.280 ;
        RECT 1201.590 43.220 1201.910 43.280 ;
      LAYER via ;
        RECT 1201.620 1678.280 1201.880 1678.540 ;
        RECT 1203.920 1678.280 1204.180 1678.540 ;
        RECT 525.880 43.220 526.140 43.480 ;
        RECT 1201.620 43.220 1201.880 43.480 ;
      LAYER met2 ;
        RECT 1203.820 1700.340 1204.100 1704.000 ;
        RECT 1203.820 1700.000 1204.120 1700.340 ;
        RECT 1203.980 1678.570 1204.120 1700.000 ;
        RECT 1201.620 1678.250 1201.880 1678.570 ;
        RECT 1203.920 1678.250 1204.180 1678.570 ;
        RECT 1201.680 43.510 1201.820 1678.250 ;
        RECT 525.880 43.190 526.140 43.510 ;
        RECT 1201.620 43.190 1201.880 43.510 ;
        RECT 525.940 2.400 526.080 43.190 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 543.790 43.080 544.110 43.140 ;
        RECT 1205.730 43.080 1206.050 43.140 ;
        RECT 543.790 42.940 1206.050 43.080 ;
        RECT 543.790 42.880 544.110 42.940 ;
        RECT 1205.730 42.880 1206.050 42.940 ;
      LAYER via ;
        RECT 543.820 42.880 544.080 43.140 ;
        RECT 1205.760 42.880 1206.020 43.140 ;
      LAYER met2 ;
        RECT 1205.660 1700.340 1205.940 1704.000 ;
        RECT 1205.660 1700.000 1205.960 1700.340 ;
        RECT 1205.820 43.170 1205.960 1700.000 ;
        RECT 543.820 42.850 544.080 43.170 ;
        RECT 1205.760 42.850 1206.020 43.170 ;
        RECT 543.880 2.400 544.020 42.850 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1207.570 1668.960 1207.890 1669.020 ;
        RECT 1209.410 1668.960 1209.730 1669.020 ;
        RECT 1207.570 1668.820 1209.730 1668.960 ;
        RECT 1207.570 1668.760 1207.890 1668.820 ;
        RECT 1209.410 1668.760 1209.730 1668.820 ;
        RECT 561.730 42.740 562.050 42.800 ;
        RECT 1209.410 42.740 1209.730 42.800 ;
        RECT 561.730 42.600 1209.730 42.740 ;
        RECT 561.730 42.540 562.050 42.600 ;
        RECT 1209.410 42.540 1209.730 42.600 ;
      LAYER via ;
        RECT 1207.600 1668.760 1207.860 1669.020 ;
        RECT 1209.440 1668.760 1209.700 1669.020 ;
        RECT 561.760 42.540 562.020 42.800 ;
        RECT 1209.440 42.540 1209.700 42.800 ;
      LAYER met2 ;
        RECT 1207.500 1700.340 1207.780 1704.000 ;
        RECT 1207.500 1700.000 1207.800 1700.340 ;
        RECT 1207.660 1669.050 1207.800 1700.000 ;
        RECT 1207.600 1668.730 1207.860 1669.050 ;
        RECT 1209.440 1668.730 1209.700 1669.050 ;
        RECT 1209.500 42.830 1209.640 1668.730 ;
        RECT 561.760 42.510 562.020 42.830 ;
        RECT 1209.440 42.510 1209.700 42.830 ;
        RECT 561.820 2.400 561.960 42.510 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 579.670 42.400 579.990 42.460 ;
        RECT 1208.950 42.400 1209.270 42.460 ;
        RECT 579.670 42.260 1209.270 42.400 ;
        RECT 579.670 42.200 579.990 42.260 ;
        RECT 1208.950 42.200 1209.270 42.260 ;
      LAYER via ;
        RECT 579.700 42.200 579.960 42.460 ;
        RECT 1208.980 42.200 1209.240 42.460 ;
      LAYER met2 ;
        RECT 1209.340 1700.410 1209.620 1704.000 ;
        RECT 1209.040 1700.270 1209.620 1700.410 ;
        RECT 1209.040 42.490 1209.180 1700.270 ;
        RECT 1209.340 1700.000 1209.620 1700.270 ;
        RECT 579.700 42.170 579.960 42.490 ;
        RECT 1208.980 42.170 1209.240 42.490 ;
        RECT 579.760 2.400 579.900 42.170 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 44.780 86.410 44.840 ;
        RECT 1158.350 44.780 1158.670 44.840 ;
        RECT 86.090 44.640 1158.670 44.780 ;
        RECT 86.090 44.580 86.410 44.640 ;
        RECT 1158.350 44.580 1158.670 44.640 ;
      LAYER via ;
        RECT 86.120 44.580 86.380 44.840 ;
        RECT 1158.380 44.580 1158.640 44.840 ;
      LAYER met2 ;
        RECT 1158.280 1700.340 1158.560 1704.000 ;
        RECT 1158.280 1700.000 1158.580 1700.340 ;
        RECT 1158.440 44.870 1158.580 1700.000 ;
        RECT 86.120 44.550 86.380 44.870 ;
        RECT 1158.380 44.550 1158.640 44.870 ;
        RECT 86.180 2.400 86.320 44.550 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 597.150 42.060 597.470 42.120 ;
        RECT 1211.250 42.060 1211.570 42.120 ;
        RECT 597.150 41.920 1211.570 42.060 ;
        RECT 597.150 41.860 597.470 41.920 ;
        RECT 1211.250 41.860 1211.570 41.920 ;
      LAYER via ;
        RECT 597.180 41.860 597.440 42.120 ;
        RECT 1211.280 41.860 1211.540 42.120 ;
      LAYER met2 ;
        RECT 1211.180 1700.340 1211.460 1704.000 ;
        RECT 1211.180 1700.000 1211.480 1700.340 ;
        RECT 1211.340 42.150 1211.480 1700.000 ;
        RECT 597.180 41.830 597.440 42.150 ;
        RECT 1211.280 41.830 1211.540 42.150 ;
        RECT 597.240 2.400 597.380 41.830 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 615.090 41.720 615.410 41.780 ;
        RECT 1213.090 41.720 1213.410 41.780 ;
        RECT 615.090 41.580 1213.410 41.720 ;
        RECT 615.090 41.520 615.410 41.580 ;
        RECT 1213.090 41.520 1213.410 41.580 ;
      LAYER via ;
        RECT 615.120 41.520 615.380 41.780 ;
        RECT 1213.120 41.520 1213.380 41.780 ;
      LAYER met2 ;
        RECT 1213.020 1700.340 1213.300 1704.000 ;
        RECT 1213.020 1700.000 1213.320 1700.340 ;
        RECT 1213.180 41.810 1213.320 1700.000 ;
        RECT 615.120 41.490 615.380 41.810 ;
        RECT 1213.120 41.490 1213.380 41.810 ;
        RECT 615.180 2.400 615.320 41.490 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 110.010 52.260 110.330 52.320 ;
        RECT 1160.650 52.260 1160.970 52.320 ;
        RECT 110.010 52.120 1160.970 52.260 ;
        RECT 110.010 52.060 110.330 52.120 ;
        RECT 1160.650 52.060 1160.970 52.120 ;
      LAYER via ;
        RECT 110.040 52.060 110.300 52.320 ;
        RECT 1160.680 52.060 1160.940 52.320 ;
      LAYER met2 ;
        RECT 1160.580 1700.340 1160.860 1704.000 ;
        RECT 1160.580 1700.000 1160.880 1700.340 ;
        RECT 1160.740 52.350 1160.880 1700.000 ;
        RECT 110.040 52.030 110.300 52.350 ;
        RECT 1160.680 52.030 1160.940 52.350 ;
        RECT 110.100 3.130 110.240 52.030 ;
        RECT 109.640 2.990 110.240 3.130 ;
        RECT 109.640 2.400 109.780 2.990 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1161.110 1678.480 1161.430 1678.540 ;
        RECT 1162.950 1678.480 1163.270 1678.540 ;
        RECT 1161.110 1678.340 1163.270 1678.480 ;
        RECT 1161.110 1678.280 1161.430 1678.340 ;
        RECT 1162.950 1678.280 1163.270 1678.340 ;
        RECT 137.610 52.600 137.930 52.660 ;
        RECT 1161.110 52.600 1161.430 52.660 ;
        RECT 137.610 52.460 1161.430 52.600 ;
        RECT 137.610 52.400 137.930 52.460 ;
        RECT 1161.110 52.400 1161.430 52.460 ;
        RECT 133.470 17.580 133.790 17.640 ;
        RECT 137.610 17.580 137.930 17.640 ;
        RECT 133.470 17.440 137.930 17.580 ;
        RECT 133.470 17.380 133.790 17.440 ;
        RECT 137.610 17.380 137.930 17.440 ;
      LAYER via ;
        RECT 1161.140 1678.280 1161.400 1678.540 ;
        RECT 1162.980 1678.280 1163.240 1678.540 ;
        RECT 137.640 52.400 137.900 52.660 ;
        RECT 1161.140 52.400 1161.400 52.660 ;
        RECT 133.500 17.380 133.760 17.640 ;
        RECT 137.640 17.380 137.900 17.640 ;
      LAYER met2 ;
        RECT 1163.340 1700.410 1163.620 1704.000 ;
        RECT 1163.040 1700.270 1163.620 1700.410 ;
        RECT 1163.040 1678.570 1163.180 1700.270 ;
        RECT 1163.340 1700.000 1163.620 1700.270 ;
        RECT 1161.140 1678.250 1161.400 1678.570 ;
        RECT 1162.980 1678.250 1163.240 1678.570 ;
        RECT 1161.200 52.690 1161.340 1678.250 ;
        RECT 137.640 52.370 137.900 52.690 ;
        RECT 1161.140 52.370 1161.400 52.690 ;
        RECT 137.700 17.670 137.840 52.370 ;
        RECT 133.500 17.350 133.760 17.670 ;
        RECT 137.640 17.350 137.900 17.670 ;
        RECT 133.560 2.400 133.700 17.350 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 52.940 151.730 53.000 ;
        RECT 1165.250 52.940 1165.570 53.000 ;
        RECT 151.410 52.800 1165.570 52.940 ;
        RECT 151.410 52.740 151.730 52.800 ;
        RECT 1165.250 52.740 1165.570 52.800 ;
      LAYER via ;
        RECT 151.440 52.740 151.700 53.000 ;
        RECT 1165.280 52.740 1165.540 53.000 ;
      LAYER met2 ;
        RECT 1165.180 1700.340 1165.460 1704.000 ;
        RECT 1165.180 1700.000 1165.480 1700.340 ;
        RECT 1165.340 53.030 1165.480 1700.000 ;
        RECT 151.440 52.710 151.700 53.030 ;
        RECT 1165.280 52.710 1165.540 53.030 ;
        RECT 151.500 2.400 151.640 52.710 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1167.090 1679.160 1167.410 1679.220 ;
        RECT 1170.770 1679.160 1171.090 1679.220 ;
        RECT 1167.090 1679.020 1171.090 1679.160 ;
        RECT 1167.090 1678.960 1167.410 1679.020 ;
        RECT 1170.770 1678.960 1171.090 1679.020 ;
        RECT 172.110 1652.640 172.430 1652.700 ;
        RECT 1170.770 1652.640 1171.090 1652.700 ;
        RECT 172.110 1652.500 1171.090 1652.640 ;
        RECT 172.110 1652.440 172.430 1652.500 ;
        RECT 1170.770 1652.440 1171.090 1652.500 ;
        RECT 169.350 17.580 169.670 17.640 ;
        RECT 172.110 17.580 172.430 17.640 ;
        RECT 169.350 17.440 172.430 17.580 ;
        RECT 169.350 17.380 169.670 17.440 ;
        RECT 172.110 17.380 172.430 17.440 ;
      LAYER via ;
        RECT 1167.120 1678.960 1167.380 1679.220 ;
        RECT 1170.800 1678.960 1171.060 1679.220 ;
        RECT 172.140 1652.440 172.400 1652.700 ;
        RECT 1170.800 1652.440 1171.060 1652.700 ;
        RECT 169.380 17.380 169.640 17.640 ;
        RECT 172.140 17.380 172.400 17.640 ;
      LAYER met2 ;
        RECT 1167.020 1700.340 1167.300 1704.000 ;
        RECT 1167.020 1700.000 1167.320 1700.340 ;
        RECT 1167.180 1679.250 1167.320 1700.000 ;
        RECT 1167.120 1678.930 1167.380 1679.250 ;
        RECT 1170.800 1678.930 1171.060 1679.250 ;
        RECT 1170.860 1652.730 1171.000 1678.930 ;
        RECT 172.140 1652.410 172.400 1652.730 ;
        RECT 1170.800 1652.410 1171.060 1652.730 ;
        RECT 172.200 17.670 172.340 1652.410 ;
        RECT 169.380 17.350 169.640 17.670 ;
        RECT 172.140 17.350 172.400 17.670 ;
        RECT 169.440 2.400 169.580 17.350 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1167.090 1678.480 1167.410 1678.540 ;
        RECT 1168.470 1678.480 1168.790 1678.540 ;
        RECT 1167.090 1678.340 1168.790 1678.480 ;
        RECT 1167.090 1678.280 1167.410 1678.340 ;
        RECT 1168.470 1678.280 1168.790 1678.340 ;
        RECT 192.810 1645.500 193.130 1645.560 ;
        RECT 1167.090 1645.500 1167.410 1645.560 ;
        RECT 192.810 1645.360 1167.410 1645.500 ;
        RECT 192.810 1645.300 193.130 1645.360 ;
        RECT 1167.090 1645.300 1167.410 1645.360 ;
        RECT 186.830 17.920 187.150 17.980 ;
        RECT 192.810 17.920 193.130 17.980 ;
        RECT 186.830 17.780 193.130 17.920 ;
        RECT 186.830 17.720 187.150 17.780 ;
        RECT 192.810 17.720 193.130 17.780 ;
      LAYER via ;
        RECT 1167.120 1678.280 1167.380 1678.540 ;
        RECT 1168.500 1678.280 1168.760 1678.540 ;
        RECT 192.840 1645.300 193.100 1645.560 ;
        RECT 1167.120 1645.300 1167.380 1645.560 ;
        RECT 186.860 17.720 187.120 17.980 ;
        RECT 192.840 17.720 193.100 17.980 ;
      LAYER met2 ;
        RECT 1168.860 1700.410 1169.140 1704.000 ;
        RECT 1168.560 1700.270 1169.140 1700.410 ;
        RECT 1168.560 1678.570 1168.700 1700.270 ;
        RECT 1168.860 1700.000 1169.140 1700.270 ;
        RECT 1167.120 1678.250 1167.380 1678.570 ;
        RECT 1168.500 1678.250 1168.760 1678.570 ;
        RECT 1167.180 1645.590 1167.320 1678.250 ;
        RECT 192.840 1645.270 193.100 1645.590 ;
        RECT 1167.120 1645.270 1167.380 1645.590 ;
        RECT 192.900 18.010 193.040 1645.270 ;
        RECT 186.860 17.690 187.120 18.010 ;
        RECT 192.840 17.690 193.100 18.010 ;
        RECT 186.920 2.400 187.060 17.690 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1166.170 1679.840 1166.490 1679.900 ;
        RECT 1170.770 1679.840 1171.090 1679.900 ;
        RECT 1166.170 1679.700 1171.090 1679.840 ;
        RECT 1166.170 1679.640 1166.490 1679.700 ;
        RECT 1170.770 1679.640 1171.090 1679.700 ;
        RECT 210.290 1624.760 210.610 1624.820 ;
        RECT 1166.630 1624.760 1166.950 1624.820 ;
        RECT 210.290 1624.620 1166.950 1624.760 ;
        RECT 210.290 1624.560 210.610 1624.620 ;
        RECT 1166.630 1624.560 1166.950 1624.620 ;
        RECT 204.770 17.580 205.090 17.640 ;
        RECT 210.290 17.580 210.610 17.640 ;
        RECT 204.770 17.440 210.610 17.580 ;
        RECT 204.770 17.380 205.090 17.440 ;
        RECT 210.290 17.380 210.610 17.440 ;
      LAYER via ;
        RECT 1166.200 1679.640 1166.460 1679.900 ;
        RECT 1170.800 1679.640 1171.060 1679.900 ;
        RECT 210.320 1624.560 210.580 1624.820 ;
        RECT 1166.660 1624.560 1166.920 1624.820 ;
        RECT 204.800 17.380 205.060 17.640 ;
        RECT 210.320 17.380 210.580 17.640 ;
      LAYER met2 ;
        RECT 1170.700 1700.340 1170.980 1704.000 ;
        RECT 1170.700 1700.000 1171.000 1700.340 ;
        RECT 1170.860 1679.930 1171.000 1700.000 ;
        RECT 1166.200 1679.610 1166.460 1679.930 ;
        RECT 1170.800 1679.610 1171.060 1679.930 ;
        RECT 1166.260 1671.170 1166.400 1679.610 ;
        RECT 1166.260 1671.030 1166.860 1671.170 ;
        RECT 1166.720 1624.850 1166.860 1671.030 ;
        RECT 210.320 1624.530 210.580 1624.850 ;
        RECT 1166.660 1624.530 1166.920 1624.850 ;
        RECT 210.380 17.670 210.520 1624.530 ;
        RECT 204.800 17.350 205.060 17.670 ;
        RECT 210.320 17.350 210.580 17.670 ;
        RECT 204.860 2.400 205.000 17.350 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 230.990 1617.960 231.310 1618.020 ;
        RECT 1172.610 1617.960 1172.930 1618.020 ;
        RECT 230.990 1617.820 1172.930 1617.960 ;
        RECT 230.990 1617.760 231.310 1617.820 ;
        RECT 1172.610 1617.760 1172.930 1617.820 ;
        RECT 222.710 18.600 223.030 18.660 ;
        RECT 230.990 18.600 231.310 18.660 ;
        RECT 222.710 18.460 231.310 18.600 ;
        RECT 222.710 18.400 223.030 18.460 ;
        RECT 230.990 18.400 231.310 18.460 ;
      LAYER via ;
        RECT 231.020 1617.760 231.280 1618.020 ;
        RECT 1172.640 1617.760 1172.900 1618.020 ;
        RECT 222.740 18.400 223.000 18.660 ;
        RECT 231.020 18.400 231.280 18.660 ;
      LAYER met2 ;
        RECT 1172.540 1700.340 1172.820 1704.000 ;
        RECT 1172.540 1700.000 1172.840 1700.340 ;
        RECT 1172.700 1618.050 1172.840 1700.000 ;
        RECT 231.020 1617.730 231.280 1618.050 ;
        RECT 1172.640 1617.730 1172.900 1618.050 ;
        RECT 231.080 18.690 231.220 1617.730 ;
        RECT 222.740 18.370 223.000 18.690 ;
        RECT 231.020 18.370 231.280 18.690 ;
        RECT 222.800 2.400 222.940 18.370 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1147.845 1642.285 1148.015 1677.135 ;
        RECT 1147.385 1553.885 1147.555 1593.835 ;
        RECT 1147.385 1497.445 1147.555 1545.555 ;
        RECT 1147.845 1352.605 1148.015 1400.715 ;
        RECT 1147.845 1256.045 1148.015 1304.155 ;
        RECT 1147.845 338.045 1148.015 386.155 ;
        RECT 1147.845 241.485 1148.015 289.595 ;
        RECT 1147.845 144.925 1148.015 193.035 ;
      LAYER mcon ;
        RECT 1147.845 1676.965 1148.015 1677.135 ;
        RECT 1147.385 1593.665 1147.555 1593.835 ;
        RECT 1147.385 1545.385 1147.555 1545.555 ;
        RECT 1147.845 1400.545 1148.015 1400.715 ;
        RECT 1147.845 1303.985 1148.015 1304.155 ;
        RECT 1147.845 385.985 1148.015 386.155 ;
        RECT 1147.845 289.425 1148.015 289.595 ;
        RECT 1147.845 192.865 1148.015 193.035 ;
      LAYER met1 ;
        RECT 1147.785 1677.120 1148.075 1677.165 ;
        RECT 1151.450 1677.120 1151.770 1677.180 ;
        RECT 1147.785 1676.980 1151.770 1677.120 ;
        RECT 1147.785 1676.935 1148.075 1676.980 ;
        RECT 1151.450 1676.920 1151.770 1676.980 ;
        RECT 1147.770 1642.440 1148.090 1642.500 ;
        RECT 1147.575 1642.300 1148.090 1642.440 ;
        RECT 1147.770 1642.240 1148.090 1642.300 ;
        RECT 1147.325 1593.820 1147.615 1593.865 ;
        RECT 1147.770 1593.820 1148.090 1593.880 ;
        RECT 1147.325 1593.680 1148.090 1593.820 ;
        RECT 1147.325 1593.635 1147.615 1593.680 ;
        RECT 1147.770 1593.620 1148.090 1593.680 ;
        RECT 1147.310 1554.040 1147.630 1554.100 ;
        RECT 1147.115 1553.900 1147.630 1554.040 ;
        RECT 1147.310 1553.840 1147.630 1553.900 ;
        RECT 1147.310 1545.540 1147.630 1545.600 ;
        RECT 1147.115 1545.400 1147.630 1545.540 ;
        RECT 1147.310 1545.340 1147.630 1545.400 ;
        RECT 1147.325 1497.600 1147.615 1497.645 ;
        RECT 1147.770 1497.600 1148.090 1497.660 ;
        RECT 1147.325 1497.460 1148.090 1497.600 ;
        RECT 1147.325 1497.415 1147.615 1497.460 ;
        RECT 1147.770 1497.400 1148.090 1497.460 ;
        RECT 1147.770 1400.700 1148.090 1400.760 ;
        RECT 1147.575 1400.560 1148.090 1400.700 ;
        RECT 1147.770 1400.500 1148.090 1400.560 ;
        RECT 1147.785 1352.760 1148.075 1352.805 ;
        RECT 1148.230 1352.760 1148.550 1352.820 ;
        RECT 1147.785 1352.620 1148.550 1352.760 ;
        RECT 1147.785 1352.575 1148.075 1352.620 ;
        RECT 1148.230 1352.560 1148.550 1352.620 ;
        RECT 1147.770 1304.140 1148.090 1304.200 ;
        RECT 1147.575 1304.000 1148.090 1304.140 ;
        RECT 1147.770 1303.940 1148.090 1304.000 ;
        RECT 1147.785 1256.200 1148.075 1256.245 ;
        RECT 1148.230 1256.200 1148.550 1256.260 ;
        RECT 1147.785 1256.060 1148.550 1256.200 ;
        RECT 1147.785 1256.015 1148.075 1256.060 ;
        RECT 1148.230 1256.000 1148.550 1256.060 ;
        RECT 1148.230 1159.300 1148.550 1159.360 ;
        RECT 1149.150 1159.300 1149.470 1159.360 ;
        RECT 1148.230 1159.160 1149.470 1159.300 ;
        RECT 1148.230 1159.100 1148.550 1159.160 ;
        RECT 1149.150 1159.100 1149.470 1159.160 ;
        RECT 1148.230 1062.740 1148.550 1062.800 ;
        RECT 1149.150 1062.740 1149.470 1062.800 ;
        RECT 1148.230 1062.600 1149.470 1062.740 ;
        RECT 1148.230 1062.540 1148.550 1062.600 ;
        RECT 1149.150 1062.540 1149.470 1062.600 ;
        RECT 1148.230 966.180 1148.550 966.240 ;
        RECT 1149.150 966.180 1149.470 966.240 ;
        RECT 1148.230 966.040 1149.470 966.180 ;
        RECT 1148.230 965.980 1148.550 966.040 ;
        RECT 1149.150 965.980 1149.470 966.040 ;
        RECT 1148.230 869.620 1148.550 869.680 ;
        RECT 1149.150 869.620 1149.470 869.680 ;
        RECT 1148.230 869.480 1149.470 869.620 ;
        RECT 1148.230 869.420 1148.550 869.480 ;
        RECT 1149.150 869.420 1149.470 869.480 ;
        RECT 1147.770 821.000 1148.090 821.060 ;
        RECT 1149.150 821.000 1149.470 821.060 ;
        RECT 1147.770 820.860 1149.470 821.000 ;
        RECT 1147.770 820.800 1148.090 820.860 ;
        RECT 1149.150 820.800 1149.470 820.860 ;
        RECT 1147.770 689.900 1148.090 690.160 ;
        RECT 1147.310 689.760 1147.630 689.820 ;
        RECT 1147.860 689.760 1148.000 689.900 ;
        RECT 1147.310 689.620 1148.000 689.760 ;
        RECT 1147.310 689.560 1147.630 689.620 ;
        RECT 1147.770 593.340 1148.090 593.600 ;
        RECT 1147.310 593.200 1147.630 593.260 ;
        RECT 1147.860 593.200 1148.000 593.340 ;
        RECT 1147.310 593.060 1148.000 593.200 ;
        RECT 1147.310 593.000 1147.630 593.060 ;
        RECT 1147.770 496.780 1148.090 497.040 ;
        RECT 1147.310 496.640 1147.630 496.700 ;
        RECT 1147.860 496.640 1148.000 496.780 ;
        RECT 1147.310 496.500 1148.000 496.640 ;
        RECT 1147.310 496.440 1147.630 496.500 ;
        RECT 1147.770 400.220 1148.090 400.480 ;
        RECT 1147.860 400.080 1148.000 400.220 ;
        RECT 1148.230 400.080 1148.550 400.140 ;
        RECT 1147.860 399.940 1148.550 400.080 ;
        RECT 1148.230 399.880 1148.550 399.940 ;
        RECT 1147.785 386.140 1148.075 386.185 ;
        RECT 1148.230 386.140 1148.550 386.200 ;
        RECT 1147.785 386.000 1148.550 386.140 ;
        RECT 1147.785 385.955 1148.075 386.000 ;
        RECT 1148.230 385.940 1148.550 386.000 ;
        RECT 1147.770 338.200 1148.090 338.260 ;
        RECT 1147.575 338.060 1148.090 338.200 ;
        RECT 1147.770 338.000 1148.090 338.060 ;
        RECT 1147.310 303.520 1147.630 303.580 ;
        RECT 1148.230 303.520 1148.550 303.580 ;
        RECT 1147.310 303.380 1148.550 303.520 ;
        RECT 1147.310 303.320 1147.630 303.380 ;
        RECT 1148.230 303.320 1148.550 303.380 ;
        RECT 1147.785 289.580 1148.075 289.625 ;
        RECT 1148.230 289.580 1148.550 289.640 ;
        RECT 1147.785 289.440 1148.550 289.580 ;
        RECT 1147.785 289.395 1148.075 289.440 ;
        RECT 1148.230 289.380 1148.550 289.440 ;
        RECT 1147.770 241.640 1148.090 241.700 ;
        RECT 1147.575 241.500 1148.090 241.640 ;
        RECT 1147.770 241.440 1148.090 241.500 ;
        RECT 1147.310 206.960 1147.630 207.020 ;
        RECT 1148.230 206.960 1148.550 207.020 ;
        RECT 1147.310 206.820 1148.550 206.960 ;
        RECT 1147.310 206.760 1147.630 206.820 ;
        RECT 1148.230 206.760 1148.550 206.820 ;
        RECT 1147.785 193.020 1148.075 193.065 ;
        RECT 1148.230 193.020 1148.550 193.080 ;
        RECT 1147.785 192.880 1148.550 193.020 ;
        RECT 1147.785 192.835 1148.075 192.880 ;
        RECT 1148.230 192.820 1148.550 192.880 ;
        RECT 1147.770 145.080 1148.090 145.140 ;
        RECT 1147.575 144.940 1148.090 145.080 ;
        RECT 1147.770 144.880 1148.090 144.940 ;
        RECT 1147.770 110.540 1148.090 110.800 ;
        RECT 1147.860 110.120 1148.000 110.540 ;
        RECT 1147.770 109.860 1148.090 110.120 ;
        RECT 19.850 51.580 20.170 51.640 ;
        RECT 1147.770 51.580 1148.090 51.640 ;
        RECT 19.850 51.440 1148.090 51.580 ;
        RECT 19.850 51.380 20.170 51.440 ;
        RECT 1147.770 51.380 1148.090 51.440 ;
      LAYER via ;
        RECT 1151.480 1676.920 1151.740 1677.180 ;
        RECT 1147.800 1642.240 1148.060 1642.500 ;
        RECT 1147.800 1593.620 1148.060 1593.880 ;
        RECT 1147.340 1553.840 1147.600 1554.100 ;
        RECT 1147.340 1545.340 1147.600 1545.600 ;
        RECT 1147.800 1497.400 1148.060 1497.660 ;
        RECT 1147.800 1400.500 1148.060 1400.760 ;
        RECT 1148.260 1352.560 1148.520 1352.820 ;
        RECT 1147.800 1303.940 1148.060 1304.200 ;
        RECT 1148.260 1256.000 1148.520 1256.260 ;
        RECT 1148.260 1159.100 1148.520 1159.360 ;
        RECT 1149.180 1159.100 1149.440 1159.360 ;
        RECT 1148.260 1062.540 1148.520 1062.800 ;
        RECT 1149.180 1062.540 1149.440 1062.800 ;
        RECT 1148.260 965.980 1148.520 966.240 ;
        RECT 1149.180 965.980 1149.440 966.240 ;
        RECT 1148.260 869.420 1148.520 869.680 ;
        RECT 1149.180 869.420 1149.440 869.680 ;
        RECT 1147.800 820.800 1148.060 821.060 ;
        RECT 1149.180 820.800 1149.440 821.060 ;
        RECT 1147.800 689.900 1148.060 690.160 ;
        RECT 1147.340 689.560 1147.600 689.820 ;
        RECT 1147.800 593.340 1148.060 593.600 ;
        RECT 1147.340 593.000 1147.600 593.260 ;
        RECT 1147.800 496.780 1148.060 497.040 ;
        RECT 1147.340 496.440 1147.600 496.700 ;
        RECT 1147.800 400.220 1148.060 400.480 ;
        RECT 1148.260 399.880 1148.520 400.140 ;
        RECT 1148.260 385.940 1148.520 386.200 ;
        RECT 1147.800 338.000 1148.060 338.260 ;
        RECT 1147.340 303.320 1147.600 303.580 ;
        RECT 1148.260 303.320 1148.520 303.580 ;
        RECT 1148.260 289.380 1148.520 289.640 ;
        RECT 1147.800 241.440 1148.060 241.700 ;
        RECT 1147.340 206.760 1147.600 207.020 ;
        RECT 1148.260 206.760 1148.520 207.020 ;
        RECT 1148.260 192.820 1148.520 193.080 ;
        RECT 1147.800 144.880 1148.060 145.140 ;
        RECT 1147.800 110.540 1148.060 110.800 ;
        RECT 1147.800 109.860 1148.060 110.120 ;
        RECT 19.880 51.380 20.140 51.640 ;
        RECT 1147.800 51.380 1148.060 51.640 ;
      LAYER met2 ;
        RECT 1151.380 1700.340 1151.660 1704.000 ;
        RECT 1151.380 1700.000 1151.680 1700.340 ;
        RECT 1151.540 1677.210 1151.680 1700.000 ;
        RECT 1151.480 1676.890 1151.740 1677.210 ;
        RECT 1147.800 1642.210 1148.060 1642.530 ;
        RECT 1147.860 1593.910 1148.000 1642.210 ;
        RECT 1147.800 1593.590 1148.060 1593.910 ;
        RECT 1147.340 1553.810 1147.600 1554.130 ;
        RECT 1147.400 1545.630 1147.540 1553.810 ;
        RECT 1147.340 1545.310 1147.600 1545.630 ;
        RECT 1147.800 1497.370 1148.060 1497.690 ;
        RECT 1147.860 1472.610 1148.000 1497.370 ;
        RECT 1147.860 1472.470 1148.460 1472.610 ;
        RECT 1148.320 1414.130 1148.460 1472.470 ;
        RECT 1147.860 1413.990 1148.460 1414.130 ;
        RECT 1147.860 1400.790 1148.000 1413.990 ;
        RECT 1147.800 1400.470 1148.060 1400.790 ;
        RECT 1148.260 1352.530 1148.520 1352.850 ;
        RECT 1148.320 1317.570 1148.460 1352.530 ;
        RECT 1147.860 1317.430 1148.460 1317.570 ;
        RECT 1147.860 1304.230 1148.000 1317.430 ;
        RECT 1147.800 1303.910 1148.060 1304.230 ;
        RECT 1148.260 1255.970 1148.520 1256.290 ;
        RECT 1148.320 1221.010 1148.460 1255.970 ;
        RECT 1147.860 1220.870 1148.460 1221.010 ;
        RECT 1147.860 1207.525 1148.000 1220.870 ;
        RECT 1147.790 1207.155 1148.070 1207.525 ;
        RECT 1149.170 1207.155 1149.450 1207.525 ;
        RECT 1149.240 1159.390 1149.380 1207.155 ;
        RECT 1148.260 1159.070 1148.520 1159.390 ;
        RECT 1149.180 1159.070 1149.440 1159.390 ;
        RECT 1148.320 1124.450 1148.460 1159.070 ;
        RECT 1147.860 1124.310 1148.460 1124.450 ;
        RECT 1147.860 1110.965 1148.000 1124.310 ;
        RECT 1147.790 1110.595 1148.070 1110.965 ;
        RECT 1149.170 1110.595 1149.450 1110.965 ;
        RECT 1149.240 1062.830 1149.380 1110.595 ;
        RECT 1148.260 1062.510 1148.520 1062.830 ;
        RECT 1149.180 1062.510 1149.440 1062.830 ;
        RECT 1148.320 1027.890 1148.460 1062.510 ;
        RECT 1147.860 1027.750 1148.460 1027.890 ;
        RECT 1147.860 1014.405 1148.000 1027.750 ;
        RECT 1147.790 1014.035 1148.070 1014.405 ;
        RECT 1149.170 1014.035 1149.450 1014.405 ;
        RECT 1149.240 966.270 1149.380 1014.035 ;
        RECT 1148.260 965.950 1148.520 966.270 ;
        RECT 1149.180 965.950 1149.440 966.270 ;
        RECT 1148.320 931.330 1148.460 965.950 ;
        RECT 1147.860 931.190 1148.460 931.330 ;
        RECT 1147.860 917.845 1148.000 931.190 ;
        RECT 1147.790 917.475 1148.070 917.845 ;
        RECT 1149.170 917.475 1149.450 917.845 ;
        RECT 1149.240 869.710 1149.380 917.475 ;
        RECT 1148.260 869.390 1148.520 869.710 ;
        RECT 1149.180 869.390 1149.440 869.710 ;
        RECT 1148.320 834.770 1148.460 869.390 ;
        RECT 1147.860 834.630 1148.460 834.770 ;
        RECT 1147.860 821.090 1148.000 834.630 ;
        RECT 1147.800 820.770 1148.060 821.090 ;
        RECT 1149.180 820.770 1149.440 821.090 ;
        RECT 1149.240 773.005 1149.380 820.770 ;
        RECT 1148.250 772.635 1148.530 773.005 ;
        RECT 1149.170 772.635 1149.450 773.005 ;
        RECT 1148.320 738.210 1148.460 772.635 ;
        RECT 1147.860 738.070 1148.460 738.210 ;
        RECT 1147.860 690.190 1148.000 738.070 ;
        RECT 1147.800 689.870 1148.060 690.190 ;
        RECT 1147.340 689.530 1147.600 689.850 ;
        RECT 1147.400 676.445 1147.540 689.530 ;
        RECT 1147.330 676.075 1147.610 676.445 ;
        RECT 1148.250 676.075 1148.530 676.445 ;
        RECT 1148.320 641.650 1148.460 676.075 ;
        RECT 1147.860 641.510 1148.460 641.650 ;
        RECT 1147.860 593.630 1148.000 641.510 ;
        RECT 1147.800 593.310 1148.060 593.630 ;
        RECT 1147.340 592.970 1147.600 593.290 ;
        RECT 1147.400 579.885 1147.540 592.970 ;
        RECT 1147.330 579.515 1147.610 579.885 ;
        RECT 1148.250 579.515 1148.530 579.885 ;
        RECT 1148.320 545.090 1148.460 579.515 ;
        RECT 1147.860 544.950 1148.460 545.090 ;
        RECT 1147.860 497.070 1148.000 544.950 ;
        RECT 1147.800 496.750 1148.060 497.070 ;
        RECT 1147.340 496.410 1147.600 496.730 ;
        RECT 1147.400 483.325 1147.540 496.410 ;
        RECT 1147.330 482.955 1147.610 483.325 ;
        RECT 1148.250 482.955 1148.530 483.325 ;
        RECT 1148.320 448.530 1148.460 482.955 ;
        RECT 1147.860 448.390 1148.460 448.530 ;
        RECT 1147.860 400.510 1148.000 448.390 ;
        RECT 1147.800 400.190 1148.060 400.510 ;
        RECT 1148.260 399.850 1148.520 400.170 ;
        RECT 1148.320 386.230 1148.460 399.850 ;
        RECT 1148.260 385.910 1148.520 386.230 ;
        RECT 1147.800 337.970 1148.060 338.290 ;
        RECT 1147.860 303.690 1148.000 337.970 ;
        RECT 1147.400 303.610 1148.000 303.690 ;
        RECT 1147.340 303.550 1148.000 303.610 ;
        RECT 1147.340 303.290 1147.600 303.550 ;
        RECT 1148.260 303.290 1148.520 303.610 ;
        RECT 1148.320 289.670 1148.460 303.290 ;
        RECT 1148.260 289.350 1148.520 289.670 ;
        RECT 1147.800 241.410 1148.060 241.730 ;
        RECT 1147.860 207.130 1148.000 241.410 ;
        RECT 1147.400 207.050 1148.000 207.130 ;
        RECT 1147.340 206.990 1148.000 207.050 ;
        RECT 1147.340 206.730 1147.600 206.990 ;
        RECT 1148.260 206.730 1148.520 207.050 ;
        RECT 1148.320 193.110 1148.460 206.730 ;
        RECT 1148.260 192.790 1148.520 193.110 ;
        RECT 1147.800 144.850 1148.060 145.170 ;
        RECT 1147.860 110.830 1148.000 144.850 ;
        RECT 1147.800 110.510 1148.060 110.830 ;
        RECT 1147.800 109.830 1148.060 110.150 ;
        RECT 1147.860 51.670 1148.000 109.830 ;
        RECT 19.880 51.350 20.140 51.670 ;
        RECT 1147.800 51.350 1148.060 51.670 ;
        RECT 19.940 3.130 20.080 51.350 ;
        RECT 19.940 2.990 20.540 3.130 ;
        RECT 20.400 2.400 20.540 2.990 ;
        RECT 20.190 -4.800 20.750 2.400 ;
      LAYER via2 ;
        RECT 1147.790 1207.200 1148.070 1207.480 ;
        RECT 1149.170 1207.200 1149.450 1207.480 ;
        RECT 1147.790 1110.640 1148.070 1110.920 ;
        RECT 1149.170 1110.640 1149.450 1110.920 ;
        RECT 1147.790 1014.080 1148.070 1014.360 ;
        RECT 1149.170 1014.080 1149.450 1014.360 ;
        RECT 1147.790 917.520 1148.070 917.800 ;
        RECT 1149.170 917.520 1149.450 917.800 ;
        RECT 1148.250 772.680 1148.530 772.960 ;
        RECT 1149.170 772.680 1149.450 772.960 ;
        RECT 1147.330 676.120 1147.610 676.400 ;
        RECT 1148.250 676.120 1148.530 676.400 ;
        RECT 1147.330 579.560 1147.610 579.840 ;
        RECT 1148.250 579.560 1148.530 579.840 ;
        RECT 1147.330 483.000 1147.610 483.280 ;
        RECT 1148.250 483.000 1148.530 483.280 ;
      LAYER met3 ;
        RECT 1147.765 1207.490 1148.095 1207.505 ;
        RECT 1149.145 1207.490 1149.475 1207.505 ;
        RECT 1147.765 1207.190 1149.475 1207.490 ;
        RECT 1147.765 1207.175 1148.095 1207.190 ;
        RECT 1149.145 1207.175 1149.475 1207.190 ;
        RECT 1147.765 1110.930 1148.095 1110.945 ;
        RECT 1149.145 1110.930 1149.475 1110.945 ;
        RECT 1147.765 1110.630 1149.475 1110.930 ;
        RECT 1147.765 1110.615 1148.095 1110.630 ;
        RECT 1149.145 1110.615 1149.475 1110.630 ;
        RECT 1147.765 1014.370 1148.095 1014.385 ;
        RECT 1149.145 1014.370 1149.475 1014.385 ;
        RECT 1147.765 1014.070 1149.475 1014.370 ;
        RECT 1147.765 1014.055 1148.095 1014.070 ;
        RECT 1149.145 1014.055 1149.475 1014.070 ;
        RECT 1147.765 917.810 1148.095 917.825 ;
        RECT 1149.145 917.810 1149.475 917.825 ;
        RECT 1147.765 917.510 1149.475 917.810 ;
        RECT 1147.765 917.495 1148.095 917.510 ;
        RECT 1149.145 917.495 1149.475 917.510 ;
        RECT 1148.225 772.970 1148.555 772.985 ;
        RECT 1149.145 772.970 1149.475 772.985 ;
        RECT 1148.225 772.670 1149.475 772.970 ;
        RECT 1148.225 772.655 1148.555 772.670 ;
        RECT 1149.145 772.655 1149.475 772.670 ;
        RECT 1147.305 676.410 1147.635 676.425 ;
        RECT 1148.225 676.410 1148.555 676.425 ;
        RECT 1147.305 676.110 1148.555 676.410 ;
        RECT 1147.305 676.095 1147.635 676.110 ;
        RECT 1148.225 676.095 1148.555 676.110 ;
        RECT 1147.305 579.850 1147.635 579.865 ;
        RECT 1148.225 579.850 1148.555 579.865 ;
        RECT 1147.305 579.550 1148.555 579.850 ;
        RECT 1147.305 579.535 1147.635 579.550 ;
        RECT 1148.225 579.535 1148.555 579.550 ;
        RECT 1147.305 483.290 1147.635 483.305 ;
        RECT 1148.225 483.290 1148.555 483.305 ;
        RECT 1147.305 482.990 1148.555 483.290 ;
        RECT 1147.305 482.975 1147.635 482.990 ;
        RECT 1148.225 482.975 1148.555 482.990 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.910 51.920 48.230 51.980 ;
        RECT 1154.210 51.920 1154.530 51.980 ;
        RECT 47.910 51.780 1154.530 51.920 ;
        RECT 47.910 51.720 48.230 51.780 ;
        RECT 1154.210 51.720 1154.530 51.780 ;
        RECT 44.230 17.580 44.550 17.640 ;
        RECT 47.910 17.580 48.230 17.640 ;
        RECT 44.230 17.440 48.230 17.580 ;
        RECT 44.230 17.380 44.550 17.440 ;
        RECT 47.910 17.380 48.230 17.440 ;
      LAYER via ;
        RECT 47.940 51.720 48.200 51.980 ;
        RECT 1154.240 51.720 1154.500 51.980 ;
        RECT 44.260 17.380 44.520 17.640 ;
        RECT 47.940 17.380 48.200 17.640 ;
      LAYER met2 ;
        RECT 1154.140 1700.340 1154.420 1704.000 ;
        RECT 1154.140 1700.000 1154.440 1700.340 ;
        RECT 1154.300 52.010 1154.440 1700.000 ;
        RECT 47.940 51.690 48.200 52.010 ;
        RECT 1154.240 51.690 1154.500 52.010 ;
        RECT 48.000 17.670 48.140 51.690 ;
        RECT 44.260 17.350 44.520 17.670 ;
        RECT 47.940 17.350 48.200 17.670 ;
        RECT 44.320 2.400 44.460 17.350 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 248.010 1659.440 248.330 1659.500 ;
        RECT 1174.910 1659.440 1175.230 1659.500 ;
        RECT 248.010 1659.300 1175.230 1659.440 ;
        RECT 248.010 1659.240 248.330 1659.300 ;
        RECT 1174.910 1659.240 1175.230 1659.300 ;
      LAYER via ;
        RECT 248.040 1659.240 248.300 1659.500 ;
        RECT 1174.940 1659.240 1175.200 1659.500 ;
      LAYER met2 ;
        RECT 1174.840 1700.340 1175.120 1704.000 ;
        RECT 1174.840 1700.000 1175.140 1700.340 ;
        RECT 1175.000 1659.530 1175.140 1700.000 ;
        RECT 248.040 1659.210 248.300 1659.530 ;
        RECT 1174.940 1659.210 1175.200 1659.530 ;
        RECT 248.100 17.410 248.240 1659.210 ;
        RECT 246.720 17.270 248.240 17.410 ;
        RECT 246.720 2.400 246.860 17.270 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 268.710 1638.700 269.030 1638.760 ;
        RECT 1176.750 1638.700 1177.070 1638.760 ;
        RECT 268.710 1638.560 1177.070 1638.700 ;
        RECT 268.710 1638.500 269.030 1638.560 ;
        RECT 1176.750 1638.500 1177.070 1638.560 ;
        RECT 264.110 17.920 264.430 17.980 ;
        RECT 268.710 17.920 269.030 17.980 ;
        RECT 264.110 17.780 269.030 17.920 ;
        RECT 264.110 17.720 264.430 17.780 ;
        RECT 268.710 17.720 269.030 17.780 ;
      LAYER via ;
        RECT 268.740 1638.500 269.000 1638.760 ;
        RECT 1176.780 1638.500 1177.040 1638.760 ;
        RECT 264.140 17.720 264.400 17.980 ;
        RECT 268.740 17.720 269.000 17.980 ;
      LAYER met2 ;
        RECT 1176.680 1700.340 1176.960 1704.000 ;
        RECT 1176.680 1700.000 1176.980 1700.340 ;
        RECT 1176.840 1638.790 1176.980 1700.000 ;
        RECT 268.740 1638.470 269.000 1638.790 ;
        RECT 1176.780 1638.470 1177.040 1638.790 ;
        RECT 268.800 18.010 268.940 1638.470 ;
        RECT 264.140 17.690 264.400 18.010 ;
        RECT 268.740 17.690 269.000 18.010 ;
        RECT 264.200 2.400 264.340 17.690 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1178.590 1656.180 1178.910 1656.440 ;
        RECT 1178.680 1655.760 1178.820 1656.180 ;
        RECT 1178.590 1655.500 1178.910 1655.760 ;
        RECT 282.050 1632.240 282.370 1632.300 ;
        RECT 1178.590 1632.240 1178.910 1632.300 ;
        RECT 282.050 1632.100 1178.910 1632.240 ;
        RECT 282.050 1632.040 282.370 1632.100 ;
        RECT 1178.590 1632.040 1178.910 1632.100 ;
      LAYER via ;
        RECT 1178.620 1656.180 1178.880 1656.440 ;
        RECT 1178.620 1655.500 1178.880 1655.760 ;
        RECT 282.080 1632.040 282.340 1632.300 ;
        RECT 1178.620 1632.040 1178.880 1632.300 ;
      LAYER met2 ;
        RECT 1178.520 1700.340 1178.800 1704.000 ;
        RECT 1178.520 1700.000 1178.820 1700.340 ;
        RECT 1178.680 1656.470 1178.820 1700.000 ;
        RECT 1178.620 1656.150 1178.880 1656.470 ;
        RECT 1178.620 1655.470 1178.880 1655.790 ;
        RECT 1178.680 1632.330 1178.820 1655.470 ;
        RECT 282.080 1632.010 282.340 1632.330 ;
        RECT 1178.620 1632.010 1178.880 1632.330 ;
        RECT 282.140 2.400 282.280 1632.010 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1180.430 1678.280 1180.750 1678.540 ;
        RECT 1180.520 1676.100 1180.660 1678.280 ;
        RECT 1184.110 1676.100 1184.430 1676.160 ;
        RECT 1180.520 1675.960 1184.430 1676.100 ;
        RECT 1184.110 1675.900 1184.430 1675.960 ;
        RECT 303.210 53.280 303.530 53.340 ;
        RECT 1184.110 53.280 1184.430 53.340 ;
        RECT 303.210 53.140 1184.430 53.280 ;
        RECT 303.210 53.080 303.530 53.140 ;
        RECT 1184.110 53.080 1184.430 53.140 ;
        RECT 299.990 16.900 300.310 16.960 ;
        RECT 303.210 16.900 303.530 16.960 ;
        RECT 299.990 16.760 303.530 16.900 ;
        RECT 299.990 16.700 300.310 16.760 ;
        RECT 303.210 16.700 303.530 16.760 ;
      LAYER via ;
        RECT 1180.460 1678.280 1180.720 1678.540 ;
        RECT 1184.140 1675.900 1184.400 1676.160 ;
        RECT 303.240 53.080 303.500 53.340 ;
        RECT 1184.140 53.080 1184.400 53.340 ;
        RECT 300.020 16.700 300.280 16.960 ;
        RECT 303.240 16.700 303.500 16.960 ;
      LAYER met2 ;
        RECT 1180.360 1700.340 1180.640 1704.000 ;
        RECT 1180.360 1700.000 1180.660 1700.340 ;
        RECT 1180.520 1678.570 1180.660 1700.000 ;
        RECT 1180.460 1678.250 1180.720 1678.570 ;
        RECT 1184.140 1675.870 1184.400 1676.190 ;
        RECT 1184.200 53.370 1184.340 1675.870 ;
        RECT 303.240 53.050 303.500 53.370 ;
        RECT 1184.140 53.050 1184.400 53.370 ;
        RECT 303.300 16.990 303.440 53.050 ;
        RECT 300.020 16.670 300.280 16.990 ;
        RECT 303.240 16.670 303.500 16.990 ;
        RECT 300.080 2.400 300.220 16.670 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 323.910 53.620 324.230 53.680 ;
        RECT 1183.650 53.620 1183.970 53.680 ;
        RECT 323.910 53.480 1183.970 53.620 ;
        RECT 323.910 53.420 324.230 53.480 ;
        RECT 1183.650 53.420 1183.970 53.480 ;
        RECT 317.930 16.900 318.250 16.960 ;
        RECT 323.910 16.900 324.230 16.960 ;
        RECT 317.930 16.760 324.230 16.900 ;
        RECT 317.930 16.700 318.250 16.760 ;
        RECT 323.910 16.700 324.230 16.760 ;
      LAYER via ;
        RECT 323.940 53.420 324.200 53.680 ;
        RECT 1183.680 53.420 1183.940 53.680 ;
        RECT 317.960 16.700 318.220 16.960 ;
        RECT 323.940 16.700 324.200 16.960 ;
      LAYER met2 ;
        RECT 1182.200 1700.340 1182.480 1704.000 ;
        RECT 1182.200 1700.000 1182.500 1700.340 ;
        RECT 1182.360 1679.840 1182.500 1700.000 ;
        RECT 1182.360 1679.700 1182.960 1679.840 ;
        RECT 1182.820 1678.650 1182.960 1679.700 ;
        RECT 1182.820 1678.510 1183.880 1678.650 ;
        RECT 1183.740 53.710 1183.880 1678.510 ;
        RECT 323.940 53.390 324.200 53.710 ;
        RECT 1183.680 53.390 1183.940 53.710 ;
        RECT 324.000 16.990 324.140 53.390 ;
        RECT 317.960 16.670 318.220 16.990 ;
        RECT 323.940 16.670 324.200 16.990 ;
        RECT 318.020 2.400 318.160 16.670 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1168.930 1683.240 1169.250 1683.300 ;
        RECT 1184.110 1683.240 1184.430 1683.300 ;
        RECT 1168.930 1683.100 1184.430 1683.240 ;
        RECT 1168.930 1683.040 1169.250 1683.100 ;
        RECT 1184.110 1683.040 1184.430 1683.100 ;
        RECT 337.710 1611.160 338.030 1611.220 ;
        RECT 1169.390 1611.160 1169.710 1611.220 ;
        RECT 337.710 1611.020 1169.710 1611.160 ;
        RECT 337.710 1610.960 338.030 1611.020 ;
        RECT 1169.390 1610.960 1169.710 1611.020 ;
      LAYER via ;
        RECT 1168.960 1683.040 1169.220 1683.300 ;
        RECT 1184.140 1683.040 1184.400 1683.300 ;
        RECT 337.740 1610.960 338.000 1611.220 ;
        RECT 1169.420 1610.960 1169.680 1611.220 ;
      LAYER met2 ;
        RECT 1184.040 1700.340 1184.320 1704.000 ;
        RECT 1184.040 1700.000 1184.340 1700.340 ;
        RECT 1184.200 1683.330 1184.340 1700.000 ;
        RECT 1168.960 1683.010 1169.220 1683.330 ;
        RECT 1184.140 1683.010 1184.400 1683.330 ;
        RECT 1169.020 1670.490 1169.160 1683.010 ;
        RECT 1169.020 1670.350 1169.620 1670.490 ;
        RECT 1169.480 1611.250 1169.620 1670.350 ;
        RECT 337.740 1610.930 338.000 1611.250 ;
        RECT 1169.420 1610.930 1169.680 1611.250 ;
        RECT 337.800 3.130 337.940 1610.930 ;
        RECT 335.960 2.990 337.940 3.130 ;
        RECT 335.960 2.400 336.100 2.990 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1185.950 1680.860 1186.270 1680.920 ;
        RECT 1179.600 1680.720 1186.270 1680.860 ;
        RECT 358.410 1680.520 358.730 1680.580 ;
        RECT 1179.600 1680.520 1179.740 1680.720 ;
        RECT 1185.950 1680.660 1186.270 1680.720 ;
        RECT 358.410 1680.380 1179.740 1680.520 ;
        RECT 358.410 1680.320 358.730 1680.380 ;
        RECT 353.350 16.900 353.670 16.960 ;
        RECT 358.410 16.900 358.730 16.960 ;
        RECT 353.350 16.760 358.730 16.900 ;
        RECT 353.350 16.700 353.670 16.760 ;
        RECT 358.410 16.700 358.730 16.760 ;
      LAYER via ;
        RECT 358.440 1680.320 358.700 1680.580 ;
        RECT 1185.980 1680.660 1186.240 1680.920 ;
        RECT 353.380 16.700 353.640 16.960 ;
        RECT 358.440 16.700 358.700 16.960 ;
      LAYER met2 ;
        RECT 1185.880 1700.340 1186.160 1704.000 ;
        RECT 1185.880 1700.000 1186.180 1700.340 ;
        RECT 1186.040 1680.950 1186.180 1700.000 ;
        RECT 1185.980 1680.630 1186.240 1680.950 ;
        RECT 358.440 1680.290 358.700 1680.610 ;
        RECT 358.500 16.990 358.640 1680.290 ;
        RECT 353.380 16.670 353.640 16.990 ;
        RECT 358.440 16.670 358.700 16.990 ;
        RECT 353.440 2.400 353.580 16.670 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.210 1673.380 372.530 1673.440 ;
        RECT 1187.790 1673.380 1188.110 1673.440 ;
        RECT 372.210 1673.240 1188.110 1673.380 ;
        RECT 372.210 1673.180 372.530 1673.240 ;
        RECT 1187.790 1673.180 1188.110 1673.240 ;
        RECT 371.290 2.960 371.610 3.020 ;
        RECT 372.210 2.960 372.530 3.020 ;
        RECT 371.290 2.820 372.530 2.960 ;
        RECT 371.290 2.760 371.610 2.820 ;
        RECT 372.210 2.760 372.530 2.820 ;
      LAYER via ;
        RECT 372.240 1673.180 372.500 1673.440 ;
        RECT 1187.820 1673.180 1188.080 1673.440 ;
        RECT 371.320 2.760 371.580 3.020 ;
        RECT 372.240 2.760 372.500 3.020 ;
      LAYER met2 ;
        RECT 1187.720 1700.340 1188.000 1704.000 ;
        RECT 1187.720 1700.000 1188.020 1700.340 ;
        RECT 1187.880 1673.470 1188.020 1700.000 ;
        RECT 372.240 1673.150 372.500 1673.470 ;
        RECT 1187.820 1673.150 1188.080 1673.470 ;
        RECT 372.300 3.050 372.440 1673.150 ;
        RECT 371.320 2.730 371.580 3.050 ;
        RECT 372.240 2.730 372.500 3.050 ;
        RECT 371.380 2.400 371.520 2.730 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 392.910 1652.980 393.230 1653.040 ;
        RECT 1189.630 1652.980 1189.950 1653.040 ;
        RECT 392.910 1652.840 1189.950 1652.980 ;
        RECT 392.910 1652.780 393.230 1652.840 ;
        RECT 1189.630 1652.780 1189.950 1652.840 ;
        RECT 389.230 16.900 389.550 16.960 ;
        RECT 392.910 16.900 393.230 16.960 ;
        RECT 389.230 16.760 393.230 16.900 ;
        RECT 389.230 16.700 389.550 16.760 ;
        RECT 392.910 16.700 393.230 16.760 ;
      LAYER via ;
        RECT 392.940 1652.780 393.200 1653.040 ;
        RECT 1189.660 1652.780 1189.920 1653.040 ;
        RECT 389.260 16.700 389.520 16.960 ;
        RECT 392.940 16.700 393.200 16.960 ;
      LAYER met2 ;
        RECT 1189.560 1700.340 1189.840 1704.000 ;
        RECT 1189.560 1700.000 1189.860 1700.340 ;
        RECT 1189.720 1653.070 1189.860 1700.000 ;
        RECT 392.940 1652.750 393.200 1653.070 ;
        RECT 1189.660 1652.750 1189.920 1653.070 ;
        RECT 393.000 16.990 393.140 1652.750 ;
        RECT 389.260 16.670 389.520 16.990 ;
        RECT 392.940 16.670 393.200 16.990 ;
        RECT 389.320 2.400 389.460 16.670 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 413.610 1604.360 413.930 1604.420 ;
        RECT 1191.470 1604.360 1191.790 1604.420 ;
        RECT 413.610 1604.220 1191.790 1604.360 ;
        RECT 413.610 1604.160 413.930 1604.220 ;
        RECT 1191.470 1604.160 1191.790 1604.220 ;
        RECT 407.170 16.900 407.490 16.960 ;
        RECT 413.610 16.900 413.930 16.960 ;
        RECT 407.170 16.760 413.930 16.900 ;
        RECT 407.170 16.700 407.490 16.760 ;
        RECT 413.610 16.700 413.930 16.760 ;
      LAYER via ;
        RECT 413.640 1604.160 413.900 1604.420 ;
        RECT 1191.500 1604.160 1191.760 1604.420 ;
        RECT 407.200 16.700 407.460 16.960 ;
        RECT 413.640 16.700 413.900 16.960 ;
      LAYER met2 ;
        RECT 1191.400 1700.340 1191.680 1704.000 ;
        RECT 1191.400 1700.000 1191.700 1700.340 ;
        RECT 1191.560 1604.450 1191.700 1700.000 ;
        RECT 413.640 1604.130 413.900 1604.450 ;
        RECT 1191.500 1604.130 1191.760 1604.450 ;
        RECT 413.700 16.990 413.840 1604.130 ;
        RECT 407.200 16.670 407.460 16.990 ;
        RECT 413.640 16.670 413.900 16.990 ;
        RECT 407.260 2.400 407.400 16.670 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1151.910 1683.920 1152.230 1683.980 ;
        RECT 1156.510 1683.920 1156.830 1683.980 ;
        RECT 1151.910 1683.780 1156.830 1683.920 ;
        RECT 1151.910 1683.720 1152.230 1683.780 ;
        RECT 1156.510 1683.720 1156.830 1683.780 ;
        RECT 68.610 1597.220 68.930 1597.280 ;
        RECT 1148.690 1597.220 1149.010 1597.280 ;
        RECT 68.610 1597.080 1149.010 1597.220 ;
        RECT 68.610 1597.020 68.930 1597.080 ;
        RECT 1148.690 1597.020 1149.010 1597.080 ;
      LAYER via ;
        RECT 1151.940 1683.720 1152.200 1683.980 ;
        RECT 1156.540 1683.720 1156.800 1683.980 ;
        RECT 68.640 1597.020 68.900 1597.280 ;
        RECT 1148.720 1597.020 1148.980 1597.280 ;
      LAYER met2 ;
        RECT 1156.440 1700.340 1156.720 1704.000 ;
        RECT 1156.440 1700.000 1156.740 1700.340 ;
        RECT 1156.600 1684.010 1156.740 1700.000 ;
        RECT 1151.940 1683.690 1152.200 1684.010 ;
        RECT 1156.540 1683.690 1156.800 1684.010 ;
        RECT 1152.000 1676.610 1152.140 1683.690 ;
        RECT 1148.780 1676.470 1152.140 1676.610 ;
        RECT 1148.780 1597.310 1148.920 1676.470 ;
        RECT 68.640 1596.990 68.900 1597.310 ;
        RECT 1148.720 1596.990 1148.980 1597.310 ;
        RECT 68.700 17.410 68.840 1596.990 ;
        RECT 68.240 17.270 68.840 17.410 ;
        RECT 68.240 2.400 68.380 17.270 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.410 1645.840 427.730 1645.900 ;
        RECT 1193.310 1645.840 1193.630 1645.900 ;
        RECT 427.410 1645.700 1193.630 1645.840 ;
        RECT 427.410 1645.640 427.730 1645.700 ;
        RECT 1193.310 1645.640 1193.630 1645.700 ;
        RECT 424.650 16.560 424.970 16.620 ;
        RECT 427.410 16.560 427.730 16.620 ;
        RECT 424.650 16.420 427.730 16.560 ;
        RECT 424.650 16.360 424.970 16.420 ;
        RECT 427.410 16.360 427.730 16.420 ;
      LAYER via ;
        RECT 427.440 1645.640 427.700 1645.900 ;
        RECT 1193.340 1645.640 1193.600 1645.900 ;
        RECT 424.680 16.360 424.940 16.620 ;
        RECT 427.440 16.360 427.700 16.620 ;
      LAYER met2 ;
        RECT 1193.240 1700.340 1193.520 1704.000 ;
        RECT 1193.240 1700.000 1193.540 1700.340 ;
        RECT 1193.400 1645.930 1193.540 1700.000 ;
        RECT 427.440 1645.610 427.700 1645.930 ;
        RECT 1193.340 1645.610 1193.600 1645.930 ;
        RECT 427.500 16.650 427.640 1645.610 ;
        RECT 424.680 16.330 424.940 16.650 ;
        RECT 427.440 16.330 427.700 16.650 ;
        RECT 424.740 2.400 424.880 16.330 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1185.490 1683.920 1185.810 1683.980 ;
        RECT 1195.150 1683.920 1195.470 1683.980 ;
        RECT 1185.490 1683.780 1195.470 1683.920 ;
        RECT 1185.490 1683.720 1185.810 1683.780 ;
        RECT 1195.150 1683.720 1195.470 1683.780 ;
        RECT 448.110 1659.780 448.430 1659.840 ;
        RECT 1185.490 1659.780 1185.810 1659.840 ;
        RECT 448.110 1659.640 1185.810 1659.780 ;
        RECT 448.110 1659.580 448.430 1659.640 ;
        RECT 1185.490 1659.580 1185.810 1659.640 ;
        RECT 442.590 15.880 442.910 15.940 ;
        RECT 448.110 15.880 448.430 15.940 ;
        RECT 442.590 15.740 448.430 15.880 ;
        RECT 442.590 15.680 442.910 15.740 ;
        RECT 448.110 15.680 448.430 15.740 ;
      LAYER via ;
        RECT 1185.520 1683.720 1185.780 1683.980 ;
        RECT 1195.180 1683.720 1195.440 1683.980 ;
        RECT 448.140 1659.580 448.400 1659.840 ;
        RECT 1185.520 1659.580 1185.780 1659.840 ;
        RECT 442.620 15.680 442.880 15.940 ;
        RECT 448.140 15.680 448.400 15.940 ;
      LAYER met2 ;
        RECT 1195.080 1700.340 1195.360 1704.000 ;
        RECT 1195.080 1700.000 1195.380 1700.340 ;
        RECT 1195.240 1684.010 1195.380 1700.000 ;
        RECT 1185.520 1683.690 1185.780 1684.010 ;
        RECT 1195.180 1683.690 1195.440 1684.010 ;
        RECT 1185.580 1659.870 1185.720 1683.690 ;
        RECT 448.140 1659.550 448.400 1659.870 ;
        RECT 1185.520 1659.550 1185.780 1659.870 ;
        RECT 448.200 15.970 448.340 1659.550 ;
        RECT 442.620 15.650 442.880 15.970 ;
        RECT 448.140 15.650 448.400 15.970 ;
        RECT 442.680 2.400 442.820 15.650 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 461.910 1666.580 462.230 1666.640 ;
        RECT 1196.990 1666.580 1197.310 1666.640 ;
        RECT 461.910 1666.440 1197.310 1666.580 ;
        RECT 461.910 1666.380 462.230 1666.440 ;
        RECT 1196.990 1666.380 1197.310 1666.440 ;
        RECT 460.530 2.960 460.850 3.020 ;
        RECT 461.910 2.960 462.230 3.020 ;
        RECT 460.530 2.820 462.230 2.960 ;
        RECT 460.530 2.760 460.850 2.820 ;
        RECT 461.910 2.760 462.230 2.820 ;
      LAYER via ;
        RECT 461.940 1666.380 462.200 1666.640 ;
        RECT 1197.020 1666.380 1197.280 1666.640 ;
        RECT 460.560 2.760 460.820 3.020 ;
        RECT 461.940 2.760 462.200 3.020 ;
      LAYER met2 ;
        RECT 1196.920 1700.340 1197.200 1704.000 ;
        RECT 1196.920 1700.000 1197.220 1700.340 ;
        RECT 1197.080 1666.670 1197.220 1700.000 ;
        RECT 461.940 1666.350 462.200 1666.670 ;
        RECT 1197.020 1666.350 1197.280 1666.670 ;
        RECT 462.000 3.050 462.140 1666.350 ;
        RECT 460.560 2.730 460.820 3.050 ;
        RECT 461.940 2.730 462.200 3.050 ;
        RECT 460.620 2.400 460.760 2.730 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 1639.040 482.930 1639.100 ;
        RECT 1198.830 1639.040 1199.150 1639.100 ;
        RECT 482.610 1638.900 1199.150 1639.040 ;
        RECT 482.610 1638.840 482.930 1638.900 ;
        RECT 1198.830 1638.840 1199.150 1638.900 ;
        RECT 478.470 15.540 478.790 15.600 ;
        RECT 482.610 15.540 482.930 15.600 ;
        RECT 478.470 15.400 482.930 15.540 ;
        RECT 478.470 15.340 478.790 15.400 ;
        RECT 482.610 15.340 482.930 15.400 ;
      LAYER via ;
        RECT 482.640 1638.840 482.900 1639.100 ;
        RECT 1198.860 1638.840 1199.120 1639.100 ;
        RECT 478.500 15.340 478.760 15.600 ;
        RECT 482.640 15.340 482.900 15.600 ;
      LAYER met2 ;
        RECT 1198.760 1700.340 1199.040 1704.000 ;
        RECT 1198.760 1700.000 1199.060 1700.340 ;
        RECT 1198.920 1639.130 1199.060 1700.000 ;
        RECT 482.640 1638.810 482.900 1639.130 ;
        RECT 1198.860 1638.810 1199.120 1639.130 ;
        RECT 482.700 15.630 482.840 1638.810 ;
        RECT 478.500 15.310 478.760 15.630 ;
        RECT 482.640 15.310 482.900 15.630 ;
        RECT 478.560 2.400 478.700 15.310 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 496.410 1590.760 496.730 1590.820 ;
        RECT 1200.670 1590.760 1200.990 1590.820 ;
        RECT 496.410 1590.620 1200.990 1590.760 ;
        RECT 496.410 1590.560 496.730 1590.620 ;
        RECT 1200.670 1590.560 1200.990 1590.620 ;
      LAYER via ;
        RECT 496.440 1590.560 496.700 1590.820 ;
        RECT 1200.700 1590.560 1200.960 1590.820 ;
      LAYER met2 ;
        RECT 1200.600 1700.340 1200.880 1704.000 ;
        RECT 1200.600 1700.000 1200.900 1700.340 ;
        RECT 1200.760 1590.850 1200.900 1700.000 ;
        RECT 496.440 1590.530 496.700 1590.850 ;
        RECT 1200.700 1590.530 1200.960 1590.850 ;
        RECT 496.500 2.400 496.640 1590.530 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1201.130 1673.040 1201.450 1673.100 ;
        RECT 1202.510 1673.040 1202.830 1673.100 ;
        RECT 1201.130 1672.900 1202.830 1673.040 ;
        RECT 1201.130 1672.840 1201.450 1672.900 ;
        RECT 1202.510 1672.840 1202.830 1672.900 ;
        RECT 517.110 1625.100 517.430 1625.160 ;
        RECT 1201.130 1625.100 1201.450 1625.160 ;
        RECT 517.110 1624.960 1201.450 1625.100 ;
        RECT 517.110 1624.900 517.430 1624.960 ;
        RECT 1201.130 1624.900 1201.450 1624.960 ;
        RECT 513.890 15.540 514.210 15.600 ;
        RECT 517.110 15.540 517.430 15.600 ;
        RECT 513.890 15.400 517.430 15.540 ;
        RECT 513.890 15.340 514.210 15.400 ;
        RECT 517.110 15.340 517.430 15.400 ;
      LAYER via ;
        RECT 1201.160 1672.840 1201.420 1673.100 ;
        RECT 1202.540 1672.840 1202.800 1673.100 ;
        RECT 517.140 1624.900 517.400 1625.160 ;
        RECT 1201.160 1624.900 1201.420 1625.160 ;
        RECT 513.920 15.340 514.180 15.600 ;
        RECT 517.140 15.340 517.400 15.600 ;
      LAYER met2 ;
        RECT 1202.440 1700.340 1202.720 1704.000 ;
        RECT 1202.440 1700.000 1202.740 1700.340 ;
        RECT 1202.600 1673.130 1202.740 1700.000 ;
        RECT 1201.160 1672.810 1201.420 1673.130 ;
        RECT 1202.540 1672.810 1202.800 1673.130 ;
        RECT 1201.220 1625.190 1201.360 1672.810 ;
        RECT 517.140 1624.870 517.400 1625.190 ;
        RECT 1201.160 1624.870 1201.420 1625.190 ;
        RECT 517.200 15.630 517.340 1624.870 ;
        RECT 513.920 15.310 514.180 15.630 ;
        RECT 517.140 15.310 517.400 15.630 ;
        RECT 513.980 2.400 514.120 15.310 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 537.350 1548.940 537.670 1549.000 ;
        RECT 1202.510 1548.940 1202.830 1549.000 ;
        RECT 537.350 1548.800 1202.830 1548.940 ;
        RECT 537.350 1548.740 537.670 1548.800 ;
        RECT 1202.510 1548.740 1202.830 1548.800 ;
        RECT 531.830 15.540 532.150 15.600 ;
        RECT 537.350 15.540 537.670 15.600 ;
        RECT 531.830 15.400 537.670 15.540 ;
        RECT 531.830 15.340 532.150 15.400 ;
        RECT 537.350 15.340 537.670 15.400 ;
      LAYER via ;
        RECT 537.380 1548.740 537.640 1549.000 ;
        RECT 1202.540 1548.740 1202.800 1549.000 ;
        RECT 531.860 15.340 532.120 15.600 ;
        RECT 537.380 15.340 537.640 15.600 ;
      LAYER met2 ;
        RECT 1204.280 1700.340 1204.560 1704.000 ;
        RECT 1204.280 1700.000 1204.580 1700.340 ;
        RECT 1204.440 1672.530 1204.580 1700.000 ;
        RECT 1202.600 1672.390 1204.580 1672.530 ;
        RECT 1202.600 1549.030 1202.740 1672.390 ;
        RECT 537.380 1548.710 537.640 1549.030 ;
        RECT 1202.540 1548.710 1202.800 1549.030 ;
        RECT 537.440 15.630 537.580 1548.710 ;
        RECT 531.860 15.310 532.120 15.630 ;
        RECT 537.380 15.310 537.640 15.630 ;
        RECT 531.920 2.400 532.060 15.310 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1203.430 1672.020 1203.750 1672.080 ;
        RECT 1206.190 1672.020 1206.510 1672.080 ;
        RECT 1203.430 1671.880 1206.510 1672.020 ;
        RECT 1203.430 1671.820 1203.750 1671.880 ;
        RECT 1206.190 1671.820 1206.510 1671.880 ;
        RECT 551.610 1583.620 551.930 1583.680 ;
        RECT 1203.430 1583.620 1203.750 1583.680 ;
        RECT 551.610 1583.480 1203.750 1583.620 ;
        RECT 551.610 1583.420 551.930 1583.480 ;
        RECT 1203.430 1583.420 1203.750 1583.480 ;
        RECT 549.770 2.960 550.090 3.020 ;
        RECT 551.610 2.960 551.930 3.020 ;
        RECT 549.770 2.820 551.930 2.960 ;
        RECT 549.770 2.760 550.090 2.820 ;
        RECT 551.610 2.760 551.930 2.820 ;
      LAYER via ;
        RECT 1203.460 1671.820 1203.720 1672.080 ;
        RECT 1206.220 1671.820 1206.480 1672.080 ;
        RECT 551.640 1583.420 551.900 1583.680 ;
        RECT 1203.460 1583.420 1203.720 1583.680 ;
        RECT 549.800 2.760 550.060 3.020 ;
        RECT 551.640 2.760 551.900 3.020 ;
      LAYER met2 ;
        RECT 1206.120 1700.340 1206.400 1704.000 ;
        RECT 1206.120 1700.000 1206.420 1700.340 ;
        RECT 1206.280 1672.110 1206.420 1700.000 ;
        RECT 1203.460 1671.790 1203.720 1672.110 ;
        RECT 1206.220 1671.790 1206.480 1672.110 ;
        RECT 1203.520 1583.710 1203.660 1671.790 ;
        RECT 551.640 1583.390 551.900 1583.710 ;
        RECT 1203.460 1583.390 1203.720 1583.710 ;
        RECT 551.700 3.050 551.840 1583.390 ;
        RECT 549.800 2.730 550.060 3.050 ;
        RECT 551.640 2.730 551.900 3.050 ;
        RECT 549.860 2.400 550.000 2.730 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1204.810 1683.920 1205.130 1683.980 ;
        RECT 1208.030 1683.920 1208.350 1683.980 ;
        RECT 1204.810 1683.780 1208.350 1683.920 ;
        RECT 1204.810 1683.720 1205.130 1683.780 ;
        RECT 1208.030 1683.720 1208.350 1683.780 ;
        RECT 572.310 1618.300 572.630 1618.360 ;
        RECT 1203.890 1618.300 1204.210 1618.360 ;
        RECT 572.310 1618.160 1204.210 1618.300 ;
        RECT 572.310 1618.100 572.630 1618.160 ;
        RECT 1203.890 1618.100 1204.210 1618.160 ;
        RECT 567.710 14.860 568.030 14.920 ;
        RECT 572.310 14.860 572.630 14.920 ;
        RECT 567.710 14.720 572.630 14.860 ;
        RECT 567.710 14.660 568.030 14.720 ;
        RECT 572.310 14.660 572.630 14.720 ;
      LAYER via ;
        RECT 1204.840 1683.720 1205.100 1683.980 ;
        RECT 1208.060 1683.720 1208.320 1683.980 ;
        RECT 572.340 1618.100 572.600 1618.360 ;
        RECT 1203.920 1618.100 1204.180 1618.360 ;
        RECT 567.740 14.660 568.000 14.920 ;
        RECT 572.340 14.660 572.600 14.920 ;
      LAYER met2 ;
        RECT 1207.960 1700.340 1208.240 1704.000 ;
        RECT 1207.960 1700.000 1208.260 1700.340 ;
        RECT 1208.120 1684.010 1208.260 1700.000 ;
        RECT 1204.840 1683.690 1205.100 1684.010 ;
        RECT 1208.060 1683.690 1208.320 1684.010 ;
        RECT 1204.900 1671.850 1205.040 1683.690 ;
        RECT 1203.980 1671.710 1205.040 1671.850 ;
        RECT 1203.980 1618.390 1204.120 1671.710 ;
        RECT 572.340 1618.070 572.600 1618.390 ;
        RECT 1203.920 1618.070 1204.180 1618.390 ;
        RECT 572.400 14.950 572.540 1618.070 ;
        RECT 567.740 14.630 568.000 14.950 ;
        RECT 572.340 14.630 572.600 14.950 ;
        RECT 567.800 2.400 567.940 14.630 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1114.190 1686.300 1114.510 1686.360 ;
        RECT 1209.870 1686.300 1210.190 1686.360 ;
        RECT 1114.190 1686.160 1210.190 1686.300 ;
        RECT 1114.190 1686.100 1114.510 1686.160 ;
        RECT 1209.870 1686.100 1210.190 1686.160 ;
        RECT 586.110 86.260 586.430 86.320 ;
        RECT 1114.190 86.260 1114.510 86.320 ;
        RECT 586.110 86.120 1114.510 86.260 ;
        RECT 586.110 86.060 586.430 86.120 ;
        RECT 1114.190 86.060 1114.510 86.120 ;
      LAYER via ;
        RECT 1114.220 1686.100 1114.480 1686.360 ;
        RECT 1209.900 1686.100 1210.160 1686.360 ;
        RECT 586.140 86.060 586.400 86.320 ;
        RECT 1114.220 86.060 1114.480 86.320 ;
      LAYER met2 ;
        RECT 1209.800 1700.340 1210.080 1704.000 ;
        RECT 1209.800 1700.000 1210.100 1700.340 ;
        RECT 1209.960 1686.390 1210.100 1700.000 ;
        RECT 1114.220 1686.070 1114.480 1686.390 ;
        RECT 1209.900 1686.070 1210.160 1686.390 ;
        RECT 1114.280 86.350 1114.420 1686.070 ;
        RECT 586.140 86.030 586.400 86.350 ;
        RECT 1114.220 86.030 1114.480 86.350 ;
        RECT 586.200 24.210 586.340 86.030 ;
        RECT 585.740 24.070 586.340 24.210 ;
        RECT 585.740 2.400 585.880 24.070 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1157.430 1663.180 1157.750 1663.240 ;
        RECT 1158.810 1663.180 1159.130 1663.240 ;
        RECT 1157.430 1663.040 1159.130 1663.180 ;
        RECT 1157.430 1662.980 1157.750 1663.040 ;
        RECT 1158.810 1662.980 1159.130 1663.040 ;
        RECT 99.890 1631.900 100.210 1631.960 ;
        RECT 1157.430 1631.900 1157.750 1631.960 ;
        RECT 99.890 1631.760 1157.750 1631.900 ;
        RECT 99.890 1631.700 100.210 1631.760 ;
        RECT 1157.430 1631.700 1157.750 1631.760 ;
        RECT 91.610 17.580 91.930 17.640 ;
        RECT 99.890 17.580 100.210 17.640 ;
        RECT 91.610 17.440 100.210 17.580 ;
        RECT 91.610 17.380 91.930 17.440 ;
        RECT 99.890 17.380 100.210 17.440 ;
      LAYER via ;
        RECT 1157.460 1662.980 1157.720 1663.240 ;
        RECT 1158.840 1662.980 1159.100 1663.240 ;
        RECT 99.920 1631.700 100.180 1631.960 ;
        RECT 1157.460 1631.700 1157.720 1631.960 ;
        RECT 91.640 17.380 91.900 17.640 ;
        RECT 99.920 17.380 100.180 17.640 ;
      LAYER met2 ;
        RECT 1158.740 1700.340 1159.020 1704.000 ;
        RECT 1158.740 1700.000 1159.040 1700.340 ;
        RECT 1158.900 1663.270 1159.040 1700.000 ;
        RECT 1157.460 1662.950 1157.720 1663.270 ;
        RECT 1158.840 1662.950 1159.100 1663.270 ;
        RECT 1157.520 1631.990 1157.660 1662.950 ;
        RECT 99.920 1631.670 100.180 1631.990 ;
        RECT 1157.460 1631.670 1157.720 1631.990 ;
        RECT 99.980 17.670 100.120 1631.670 ;
        RECT 91.640 17.350 91.900 17.670 ;
        RECT 99.920 17.350 100.180 17.670 ;
        RECT 91.700 2.400 91.840 17.350 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.810 1611.500 607.130 1611.560 ;
        RECT 1211.710 1611.500 1212.030 1611.560 ;
        RECT 606.810 1611.360 1212.030 1611.500 ;
        RECT 606.810 1611.300 607.130 1611.360 ;
        RECT 1211.710 1611.300 1212.030 1611.360 ;
        RECT 603.130 14.520 603.450 14.580 ;
        RECT 606.810 14.520 607.130 14.580 ;
        RECT 603.130 14.380 607.130 14.520 ;
        RECT 603.130 14.320 603.450 14.380 ;
        RECT 606.810 14.320 607.130 14.380 ;
      LAYER via ;
        RECT 606.840 1611.300 607.100 1611.560 ;
        RECT 1211.740 1611.300 1212.000 1611.560 ;
        RECT 603.160 14.320 603.420 14.580 ;
        RECT 606.840 14.320 607.100 14.580 ;
      LAYER met2 ;
        RECT 1211.640 1700.340 1211.920 1704.000 ;
        RECT 1211.640 1700.000 1211.940 1700.340 ;
        RECT 1211.800 1611.590 1211.940 1700.000 ;
        RECT 606.840 1611.270 607.100 1611.590 ;
        RECT 1211.740 1611.270 1212.000 1611.590 ;
        RECT 606.900 14.610 607.040 1611.270 ;
        RECT 603.160 14.290 603.420 14.610 ;
        RECT 606.840 14.290 607.100 14.610 ;
        RECT 603.220 2.400 603.360 14.290 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1212.630 1678.140 1212.950 1678.200 ;
        RECT 1213.550 1678.140 1213.870 1678.200 ;
        RECT 1212.630 1678.000 1213.870 1678.140 ;
        RECT 1212.630 1677.940 1212.950 1678.000 ;
        RECT 1213.550 1677.940 1213.870 1678.000 ;
        RECT 627.050 1604.700 627.370 1604.760 ;
        RECT 1212.630 1604.700 1212.950 1604.760 ;
        RECT 627.050 1604.560 1212.950 1604.700 ;
        RECT 627.050 1604.500 627.370 1604.560 ;
        RECT 1212.630 1604.500 1212.950 1604.560 ;
        RECT 621.070 20.980 621.390 21.040 ;
        RECT 627.050 20.980 627.370 21.040 ;
        RECT 621.070 20.840 627.370 20.980 ;
        RECT 621.070 20.780 621.390 20.840 ;
        RECT 627.050 20.780 627.370 20.840 ;
      LAYER via ;
        RECT 1212.660 1677.940 1212.920 1678.200 ;
        RECT 1213.580 1677.940 1213.840 1678.200 ;
        RECT 627.080 1604.500 627.340 1604.760 ;
        RECT 1212.660 1604.500 1212.920 1604.760 ;
        RECT 621.100 20.780 621.360 21.040 ;
        RECT 627.080 20.780 627.340 21.040 ;
      LAYER met2 ;
        RECT 1213.480 1700.340 1213.760 1704.000 ;
        RECT 1213.480 1700.000 1213.780 1700.340 ;
        RECT 1213.640 1678.230 1213.780 1700.000 ;
        RECT 1212.660 1677.910 1212.920 1678.230 ;
        RECT 1213.580 1677.910 1213.840 1678.230 ;
        RECT 1212.720 1604.790 1212.860 1677.910 ;
        RECT 627.080 1604.470 627.340 1604.790 ;
        RECT 1212.660 1604.470 1212.920 1604.790 ;
        RECT 627.140 21.070 627.280 1604.470 ;
        RECT 621.100 20.750 621.360 21.070 ;
        RECT 627.080 20.750 627.340 21.070 ;
        RECT 621.160 2.400 621.300 20.750 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1161.110 1679.500 1161.430 1679.560 ;
        RECT 1163.410 1679.500 1163.730 1679.560 ;
        RECT 1161.110 1679.360 1163.730 1679.500 ;
        RECT 1161.110 1679.300 1161.430 1679.360 ;
        RECT 1163.410 1679.300 1163.730 1679.360 ;
        RECT 120.590 1576.480 120.910 1576.540 ;
        RECT 1163.410 1576.480 1163.730 1576.540 ;
        RECT 120.590 1576.340 1163.730 1576.480 ;
        RECT 120.590 1576.280 120.910 1576.340 ;
        RECT 1163.410 1576.280 1163.730 1576.340 ;
        RECT 115.530 17.580 115.850 17.640 ;
        RECT 120.590 17.580 120.910 17.640 ;
        RECT 115.530 17.440 120.910 17.580 ;
        RECT 115.530 17.380 115.850 17.440 ;
        RECT 120.590 17.380 120.910 17.440 ;
      LAYER via ;
        RECT 1161.140 1679.300 1161.400 1679.560 ;
        RECT 1163.440 1679.300 1163.700 1679.560 ;
        RECT 120.620 1576.280 120.880 1576.540 ;
        RECT 1163.440 1576.280 1163.700 1576.540 ;
        RECT 115.560 17.380 115.820 17.640 ;
        RECT 120.620 17.380 120.880 17.640 ;
      LAYER met2 ;
        RECT 1161.500 1700.410 1161.780 1704.000 ;
        RECT 1161.200 1700.270 1161.780 1700.410 ;
        RECT 1161.200 1679.590 1161.340 1700.270 ;
        RECT 1161.500 1700.000 1161.780 1700.270 ;
        RECT 1161.140 1679.270 1161.400 1679.590 ;
        RECT 1163.440 1679.270 1163.700 1679.590 ;
        RECT 1163.500 1576.570 1163.640 1679.270 ;
        RECT 120.620 1576.250 120.880 1576.570 ;
        RECT 1163.440 1576.250 1163.700 1576.570 ;
        RECT 120.680 17.670 120.820 1576.250 ;
        RECT 115.560 17.350 115.820 17.670 ;
        RECT 120.620 17.350 120.880 17.670 ;
        RECT 115.620 2.400 115.760 17.350 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1160.190 1679.160 1160.510 1679.220 ;
        RECT 1163.870 1679.160 1164.190 1679.220 ;
        RECT 1160.190 1679.020 1164.190 1679.160 ;
        RECT 1160.190 1678.960 1160.510 1679.020 ;
        RECT 1163.870 1678.960 1164.190 1679.020 ;
        RECT 155.090 1569.680 155.410 1569.740 ;
        RECT 1160.190 1569.680 1160.510 1569.740 ;
        RECT 155.090 1569.540 1160.510 1569.680 ;
        RECT 155.090 1569.480 155.410 1569.540 ;
        RECT 1160.190 1569.480 1160.510 1569.540 ;
        RECT 139.450 16.220 139.770 16.280 ;
        RECT 155.090 16.220 155.410 16.280 ;
        RECT 139.450 16.080 155.410 16.220 ;
        RECT 139.450 16.020 139.770 16.080 ;
        RECT 155.090 16.020 155.410 16.080 ;
      LAYER via ;
        RECT 1160.220 1678.960 1160.480 1679.220 ;
        RECT 1163.900 1678.960 1164.160 1679.220 ;
        RECT 155.120 1569.480 155.380 1569.740 ;
        RECT 1160.220 1569.480 1160.480 1569.740 ;
        RECT 139.480 16.020 139.740 16.280 ;
        RECT 155.120 16.020 155.380 16.280 ;
      LAYER met2 ;
        RECT 1163.800 1700.340 1164.080 1704.000 ;
        RECT 1163.800 1700.000 1164.100 1700.340 ;
        RECT 1163.960 1679.250 1164.100 1700.000 ;
        RECT 1160.220 1678.930 1160.480 1679.250 ;
        RECT 1163.900 1678.930 1164.160 1679.250 ;
        RECT 1160.280 1569.770 1160.420 1678.930 ;
        RECT 155.120 1569.450 155.380 1569.770 ;
        RECT 1160.220 1569.450 1160.480 1569.770 ;
        RECT 155.180 16.310 155.320 1569.450 ;
        RECT 139.480 15.990 139.740 16.310 ;
        RECT 155.120 15.990 155.380 16.310 ;
        RECT 139.540 2.400 139.680 15.990 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.310 1562.880 158.630 1562.940 ;
        RECT 1165.710 1562.880 1166.030 1562.940 ;
        RECT 158.310 1562.740 1166.030 1562.880 ;
        RECT 158.310 1562.680 158.630 1562.740 ;
        RECT 1165.710 1562.680 1166.030 1562.740 ;
      LAYER via ;
        RECT 158.340 1562.680 158.600 1562.940 ;
        RECT 1165.740 1562.680 1166.000 1562.940 ;
      LAYER met2 ;
        RECT 1165.640 1700.340 1165.920 1704.000 ;
        RECT 1165.640 1700.000 1165.940 1700.340 ;
        RECT 1165.800 1562.970 1165.940 1700.000 ;
        RECT 158.340 1562.650 158.600 1562.970 ;
        RECT 1165.740 1562.650 1166.000 1562.970 ;
        RECT 158.400 17.410 158.540 1562.650 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1167.550 1656.040 1167.870 1656.100 ;
        RECT 1168.470 1656.040 1168.790 1656.100 ;
        RECT 1167.550 1655.900 1168.790 1656.040 ;
        RECT 1167.550 1655.840 1167.870 1655.900 ;
        RECT 1168.470 1655.840 1168.790 1655.900 ;
        RECT 1167.550 1608.100 1167.870 1608.160 ;
        RECT 1168.470 1608.100 1168.790 1608.160 ;
        RECT 1167.550 1607.960 1168.790 1608.100 ;
        RECT 1167.550 1607.900 1167.870 1607.960 ;
        RECT 1168.470 1607.900 1168.790 1607.960 ;
        RECT 217.190 1535.340 217.510 1535.400 ;
        RECT 1168.470 1535.340 1168.790 1535.400 ;
        RECT 217.190 1535.200 1168.790 1535.340 ;
        RECT 217.190 1535.140 217.510 1535.200 ;
        RECT 1168.470 1535.140 1168.790 1535.200 ;
        RECT 174.870 17.920 175.190 17.980 ;
        RECT 217.190 17.920 217.510 17.980 ;
        RECT 174.870 17.780 186.600 17.920 ;
        RECT 174.870 17.720 175.190 17.780 ;
        RECT 186.460 17.580 186.600 17.780 ;
        RECT 193.360 17.780 217.510 17.920 ;
        RECT 193.360 17.580 193.500 17.780 ;
        RECT 217.190 17.720 217.510 17.780 ;
        RECT 186.460 17.440 193.500 17.580 ;
      LAYER via ;
        RECT 1167.580 1655.840 1167.840 1656.100 ;
        RECT 1168.500 1655.840 1168.760 1656.100 ;
        RECT 1167.580 1607.900 1167.840 1608.160 ;
        RECT 1168.500 1607.900 1168.760 1608.160 ;
        RECT 217.220 1535.140 217.480 1535.400 ;
        RECT 1168.500 1535.140 1168.760 1535.400 ;
        RECT 174.900 17.720 175.160 17.980 ;
        RECT 217.220 17.720 217.480 17.980 ;
      LAYER met2 ;
        RECT 1167.480 1700.340 1167.760 1704.000 ;
        RECT 1167.480 1700.000 1167.780 1700.340 ;
        RECT 1167.640 1669.810 1167.780 1700.000 ;
        RECT 1167.640 1669.670 1168.700 1669.810 ;
        RECT 1168.560 1656.130 1168.700 1669.670 ;
        RECT 1167.580 1655.810 1167.840 1656.130 ;
        RECT 1168.500 1655.810 1168.760 1656.130 ;
        RECT 1167.640 1608.190 1167.780 1655.810 ;
        RECT 1167.580 1607.870 1167.840 1608.190 ;
        RECT 1168.500 1607.870 1168.760 1608.190 ;
        RECT 1168.560 1535.430 1168.700 1607.870 ;
        RECT 217.220 1535.110 217.480 1535.430 ;
        RECT 1168.500 1535.110 1168.760 1535.430 ;
        RECT 217.280 18.010 217.420 1535.110 ;
        RECT 174.900 17.690 175.160 18.010 ;
        RECT 217.220 17.690 217.480 18.010 ;
        RECT 174.960 2.400 175.100 17.690 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1168.010 1669.300 1168.330 1669.360 ;
        RECT 1170.310 1669.300 1170.630 1669.360 ;
        RECT 1168.010 1669.160 1170.630 1669.300 ;
        RECT 1168.010 1669.100 1168.330 1669.160 ;
        RECT 1170.310 1669.100 1170.630 1669.160 ;
        RECT 192.350 1528.200 192.670 1528.260 ;
        RECT 1168.010 1528.200 1168.330 1528.260 ;
        RECT 192.350 1528.060 1168.330 1528.200 ;
        RECT 192.350 1528.000 192.670 1528.060 ;
        RECT 1168.010 1528.000 1168.330 1528.060 ;
      LAYER via ;
        RECT 1168.040 1669.100 1168.300 1669.360 ;
        RECT 1170.340 1669.100 1170.600 1669.360 ;
        RECT 192.380 1528.000 192.640 1528.260 ;
        RECT 1168.040 1528.000 1168.300 1528.260 ;
      LAYER met2 ;
        RECT 1169.320 1700.340 1169.600 1704.000 ;
        RECT 1169.320 1700.000 1169.620 1700.340 ;
        RECT 1169.480 1672.530 1169.620 1700.000 ;
        RECT 1169.480 1672.390 1170.540 1672.530 ;
        RECT 1170.400 1669.390 1170.540 1672.390 ;
        RECT 1168.040 1669.070 1168.300 1669.390 ;
        RECT 1170.340 1669.070 1170.600 1669.390 ;
        RECT 1168.100 1528.290 1168.240 1669.070 ;
        RECT 192.380 1527.970 192.640 1528.290 ;
        RECT 1168.040 1527.970 1168.300 1528.290 ;
        RECT 192.440 17.410 192.580 1527.970 ;
        RECT 192.440 17.270 193.040 17.410 ;
        RECT 192.900 2.400 193.040 17.270 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 213.510 1521.400 213.830 1521.460 ;
        RECT 1171.230 1521.400 1171.550 1521.460 ;
        RECT 213.510 1521.260 1171.550 1521.400 ;
        RECT 213.510 1521.200 213.830 1521.260 ;
        RECT 1171.230 1521.200 1171.550 1521.260 ;
        RECT 210.750 17.580 211.070 17.640 ;
        RECT 213.510 17.580 213.830 17.640 ;
        RECT 210.750 17.440 213.830 17.580 ;
        RECT 210.750 17.380 211.070 17.440 ;
        RECT 213.510 17.380 213.830 17.440 ;
      LAYER via ;
        RECT 213.540 1521.200 213.800 1521.460 ;
        RECT 1171.260 1521.200 1171.520 1521.460 ;
        RECT 210.780 17.380 211.040 17.640 ;
        RECT 213.540 17.380 213.800 17.640 ;
      LAYER met2 ;
        RECT 1171.160 1700.340 1171.440 1704.000 ;
        RECT 1171.160 1700.000 1171.460 1700.340 ;
        RECT 1171.320 1521.490 1171.460 1700.000 ;
        RECT 213.540 1521.170 213.800 1521.490 ;
        RECT 1171.260 1521.170 1171.520 1521.490 ;
        RECT 213.600 17.670 213.740 1521.170 ;
        RECT 210.780 17.350 211.040 17.670 ;
        RECT 213.540 17.350 213.800 17.670 ;
        RECT 210.840 2.400 210.980 17.350 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1173.070 1678.140 1173.390 1678.200 ;
        RECT 1179.510 1678.140 1179.830 1678.200 ;
        RECT 1173.070 1678.000 1179.830 1678.140 ;
        RECT 1173.070 1677.940 1173.390 1678.000 ;
        RECT 1179.510 1677.940 1179.830 1678.000 ;
        RECT 251.690 1555.740 252.010 1555.800 ;
        RECT 1179.510 1555.740 1179.830 1555.800 ;
        RECT 251.690 1555.600 1179.830 1555.740 ;
        RECT 251.690 1555.540 252.010 1555.600 ;
        RECT 1179.510 1555.540 1179.830 1555.600 ;
        RECT 228.690 14.520 229.010 14.580 ;
        RECT 251.690 14.520 252.010 14.580 ;
        RECT 228.690 14.380 252.010 14.520 ;
        RECT 228.690 14.320 229.010 14.380 ;
        RECT 251.690 14.320 252.010 14.380 ;
      LAYER via ;
        RECT 1173.100 1677.940 1173.360 1678.200 ;
        RECT 1179.540 1677.940 1179.800 1678.200 ;
        RECT 251.720 1555.540 251.980 1555.800 ;
        RECT 1179.540 1555.540 1179.800 1555.800 ;
        RECT 228.720 14.320 228.980 14.580 ;
        RECT 251.720 14.320 251.980 14.580 ;
      LAYER met2 ;
        RECT 1173.000 1700.340 1173.280 1704.000 ;
        RECT 1173.000 1700.000 1173.300 1700.340 ;
        RECT 1173.160 1678.230 1173.300 1700.000 ;
        RECT 1173.100 1677.910 1173.360 1678.230 ;
        RECT 1179.540 1677.910 1179.800 1678.230 ;
        RECT 1179.600 1555.830 1179.740 1677.910 ;
        RECT 251.720 1555.510 251.980 1555.830 ;
        RECT 1179.540 1555.510 1179.800 1555.830 ;
        RECT 251.780 14.610 251.920 1555.510 ;
        RECT 228.720 14.290 228.980 14.610 ;
        RECT 251.720 14.290 251.980 14.610 ;
        RECT 228.780 2.400 228.920 14.290 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 72.290 1687.660 72.610 1687.720 ;
        RECT 1154.670 1687.660 1154.990 1687.720 ;
        RECT 72.290 1687.520 1154.990 1687.660 ;
        RECT 72.290 1687.460 72.610 1687.520 ;
        RECT 1154.670 1687.460 1154.990 1687.520 ;
        RECT 50.210 17.580 50.530 17.640 ;
        RECT 72.290 17.580 72.610 17.640 ;
        RECT 50.210 17.440 72.610 17.580 ;
        RECT 50.210 17.380 50.530 17.440 ;
        RECT 72.290 17.380 72.610 17.440 ;
      LAYER via ;
        RECT 72.320 1687.460 72.580 1687.720 ;
        RECT 1154.700 1687.460 1154.960 1687.720 ;
        RECT 50.240 17.380 50.500 17.640 ;
        RECT 72.320 17.380 72.580 17.640 ;
      LAYER met2 ;
        RECT 1154.600 1700.340 1154.880 1704.000 ;
        RECT 1154.600 1700.000 1154.900 1700.340 ;
        RECT 1154.760 1687.750 1154.900 1700.000 ;
        RECT 72.320 1687.430 72.580 1687.750 ;
        RECT 1154.700 1687.430 1154.960 1687.750 ;
        RECT 72.380 17.670 72.520 1687.430 ;
        RECT 50.240 17.350 50.500 17.670 ;
        RECT 72.320 17.350 72.580 17.670 ;
        RECT 50.300 2.400 50.440 17.350 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 254.910 1590.420 255.230 1590.480 ;
        RECT 1174.450 1590.420 1174.770 1590.480 ;
        RECT 254.910 1590.280 1174.770 1590.420 ;
        RECT 254.910 1590.220 255.230 1590.280 ;
        RECT 1174.450 1590.220 1174.770 1590.280 ;
        RECT 252.610 17.920 252.930 17.980 ;
        RECT 254.910 17.920 255.230 17.980 ;
        RECT 252.610 17.780 255.230 17.920 ;
        RECT 252.610 17.720 252.930 17.780 ;
        RECT 254.910 17.720 255.230 17.780 ;
      LAYER via ;
        RECT 254.940 1590.220 255.200 1590.480 ;
        RECT 1174.480 1590.220 1174.740 1590.480 ;
        RECT 252.640 17.720 252.900 17.980 ;
        RECT 254.940 17.720 255.200 17.980 ;
      LAYER met2 ;
        RECT 1175.300 1700.340 1175.580 1704.000 ;
        RECT 1175.300 1700.000 1175.600 1700.340 ;
        RECT 1175.460 1658.930 1175.600 1700.000 ;
        RECT 1174.540 1658.790 1175.600 1658.930 ;
        RECT 1174.540 1590.510 1174.680 1658.790 ;
        RECT 254.940 1590.190 255.200 1590.510 ;
        RECT 1174.480 1590.190 1174.740 1590.510 ;
        RECT 255.000 18.010 255.140 1590.190 ;
        RECT 252.640 17.690 252.900 18.010 ;
        RECT 254.940 17.690 255.200 18.010 ;
        RECT 252.700 2.400 252.840 17.690 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1176.365 1509.685 1176.535 1587.035 ;
        RECT 1176.825 1448.825 1176.995 1490.475 ;
        RECT 1175.905 1304.325 1176.075 1369.775 ;
        RECT 1175.905 1220.005 1176.075 1297.015 ;
        RECT 1175.905 786.845 1176.075 813.875 ;
        RECT 1176.365 669.545 1176.535 717.655 ;
        RECT 1176.365 614.125 1176.535 621.095 ;
        RECT 1176.365 379.525 1176.535 427.635 ;
        RECT 1175.905 186.405 1176.075 234.515 ;
      LAYER mcon ;
        RECT 1176.365 1586.865 1176.535 1587.035 ;
        RECT 1176.825 1490.305 1176.995 1490.475 ;
        RECT 1175.905 1369.605 1176.075 1369.775 ;
        RECT 1175.905 1296.845 1176.075 1297.015 ;
        RECT 1175.905 813.705 1176.075 813.875 ;
        RECT 1176.365 717.485 1176.535 717.655 ;
        RECT 1176.365 620.925 1176.535 621.095 ;
        RECT 1176.365 427.465 1176.535 427.635 ;
        RECT 1175.905 234.345 1176.075 234.515 ;
      LAYER met1 ;
        RECT 1175.830 1587.020 1176.150 1587.080 ;
        RECT 1176.305 1587.020 1176.595 1587.065 ;
        RECT 1175.830 1586.880 1176.595 1587.020 ;
        RECT 1175.830 1586.820 1176.150 1586.880 ;
        RECT 1176.305 1586.835 1176.595 1586.880 ;
        RECT 1176.305 1509.840 1176.595 1509.885 ;
        RECT 1176.750 1509.840 1177.070 1509.900 ;
        RECT 1176.305 1509.700 1177.070 1509.840 ;
        RECT 1176.305 1509.655 1176.595 1509.700 ;
        RECT 1176.750 1509.640 1177.070 1509.700 ;
        RECT 1176.750 1490.460 1177.070 1490.520 ;
        RECT 1176.555 1490.320 1177.070 1490.460 ;
        RECT 1176.750 1490.260 1177.070 1490.320 ;
        RECT 1176.750 1448.980 1177.070 1449.040 ;
        RECT 1176.555 1448.840 1177.070 1448.980 ;
        RECT 1176.750 1448.780 1177.070 1448.840 ;
        RECT 1175.830 1393.900 1176.150 1393.960 ;
        RECT 1176.750 1393.900 1177.070 1393.960 ;
        RECT 1175.830 1393.760 1177.070 1393.900 ;
        RECT 1175.830 1393.700 1176.150 1393.760 ;
        RECT 1176.750 1393.700 1177.070 1393.760 ;
        RECT 1175.845 1369.760 1176.135 1369.805 ;
        RECT 1176.290 1369.760 1176.610 1369.820 ;
        RECT 1175.845 1369.620 1176.610 1369.760 ;
        RECT 1175.845 1369.575 1176.135 1369.620 ;
        RECT 1176.290 1369.560 1176.610 1369.620 ;
        RECT 1175.830 1304.480 1176.150 1304.540 ;
        RECT 1175.635 1304.340 1176.150 1304.480 ;
        RECT 1175.830 1304.280 1176.150 1304.340 ;
        RECT 1175.830 1297.000 1176.150 1297.060 ;
        RECT 1175.635 1296.860 1176.150 1297.000 ;
        RECT 1175.830 1296.800 1176.150 1296.860 ;
        RECT 1175.830 1220.160 1176.150 1220.220 ;
        RECT 1175.635 1220.020 1176.150 1220.160 ;
        RECT 1175.830 1219.960 1176.150 1220.020 ;
        RECT 1174.910 1159.300 1175.230 1159.360 ;
        RECT 1176.290 1159.300 1176.610 1159.360 ;
        RECT 1174.910 1159.160 1176.610 1159.300 ;
        RECT 1174.910 1159.100 1175.230 1159.160 ;
        RECT 1176.290 1159.100 1176.610 1159.160 ;
        RECT 1175.830 1111.020 1176.150 1111.080 ;
        RECT 1176.750 1111.020 1177.070 1111.080 ;
        RECT 1175.830 1110.880 1177.070 1111.020 ;
        RECT 1175.830 1110.820 1176.150 1110.880 ;
        RECT 1176.750 1110.820 1177.070 1110.880 ;
        RECT 1175.830 1014.120 1176.150 1014.180 ;
        RECT 1176.290 1014.120 1176.610 1014.180 ;
        RECT 1175.830 1013.980 1176.610 1014.120 ;
        RECT 1175.830 1013.920 1176.150 1013.980 ;
        RECT 1176.290 1013.920 1176.610 1013.980 ;
        RECT 1176.290 1007.120 1176.610 1007.380 ;
        RECT 1174.910 1006.980 1175.230 1007.040 ;
        RECT 1176.380 1006.980 1176.520 1007.120 ;
        RECT 1174.910 1006.840 1176.520 1006.980 ;
        RECT 1174.910 1006.780 1175.230 1006.840 ;
        RECT 1174.910 917.900 1175.230 917.960 ;
        RECT 1175.830 917.900 1176.150 917.960 ;
        RECT 1174.910 917.760 1176.150 917.900 ;
        RECT 1174.910 917.700 1175.230 917.760 ;
        RECT 1175.830 917.700 1176.150 917.760 ;
        RECT 1174.910 869.620 1175.230 869.680 ;
        RECT 1176.290 869.620 1176.610 869.680 ;
        RECT 1174.910 869.480 1176.610 869.620 ;
        RECT 1174.910 869.420 1175.230 869.480 ;
        RECT 1176.290 869.420 1176.610 869.480 ;
        RECT 1174.910 862.480 1175.230 862.540 ;
        RECT 1176.290 862.480 1176.610 862.540 ;
        RECT 1174.910 862.340 1176.610 862.480 ;
        RECT 1174.910 862.280 1175.230 862.340 ;
        RECT 1176.290 862.280 1176.610 862.340 ;
        RECT 1175.830 813.860 1176.150 813.920 ;
        RECT 1175.635 813.720 1176.150 813.860 ;
        RECT 1175.830 813.660 1176.150 813.720 ;
        RECT 1175.830 787.000 1176.150 787.060 ;
        RECT 1175.635 786.860 1176.150 787.000 ;
        RECT 1175.830 786.800 1176.150 786.860 ;
        RECT 1175.830 724.240 1176.150 724.500 ;
        RECT 1175.920 724.100 1176.060 724.240 ;
        RECT 1176.290 724.100 1176.610 724.160 ;
        RECT 1175.920 723.960 1176.610 724.100 ;
        RECT 1176.290 723.900 1176.610 723.960 ;
        RECT 1176.290 717.640 1176.610 717.700 ;
        RECT 1176.095 717.500 1176.610 717.640 ;
        RECT 1176.290 717.440 1176.610 717.500 ;
        RECT 1176.290 669.700 1176.610 669.760 ;
        RECT 1176.095 669.560 1176.610 669.700 ;
        RECT 1176.290 669.500 1176.610 669.560 ;
        RECT 1176.290 621.080 1176.610 621.140 ;
        RECT 1176.095 620.940 1176.610 621.080 ;
        RECT 1176.290 620.880 1176.610 620.940 ;
        RECT 1176.290 614.280 1176.610 614.340 ;
        RECT 1176.095 614.140 1176.610 614.280 ;
        RECT 1176.290 614.080 1176.610 614.140 ;
        RECT 1176.290 572.460 1176.610 572.520 ;
        RECT 1176.750 572.460 1177.070 572.520 ;
        RECT 1176.290 572.320 1177.070 572.460 ;
        RECT 1176.290 572.260 1176.610 572.320 ;
        RECT 1176.750 572.260 1177.070 572.320 ;
        RECT 1176.750 497.660 1177.070 497.720 ;
        RECT 1175.920 497.520 1177.070 497.660 ;
        RECT 1175.920 497.040 1176.060 497.520 ;
        RECT 1176.750 497.460 1177.070 497.520 ;
        RECT 1175.830 496.780 1176.150 497.040 ;
        RECT 1175.830 434.760 1176.150 434.820 ;
        RECT 1176.290 434.760 1176.610 434.820 ;
        RECT 1175.830 434.620 1176.610 434.760 ;
        RECT 1175.830 434.560 1176.150 434.620 ;
        RECT 1176.290 434.560 1176.610 434.620 ;
        RECT 1176.290 427.620 1176.610 427.680 ;
        RECT 1176.095 427.480 1176.610 427.620 ;
        RECT 1176.290 427.420 1176.610 427.480 ;
        RECT 1176.290 379.680 1176.610 379.740 ;
        RECT 1176.095 379.540 1176.610 379.680 ;
        RECT 1176.290 379.480 1176.610 379.540 ;
        RECT 1176.290 352.480 1176.610 352.540 ;
        RECT 1175.920 352.340 1176.610 352.480 ;
        RECT 1175.920 351.860 1176.060 352.340 ;
        RECT 1176.290 352.280 1176.610 352.340 ;
        RECT 1175.830 351.600 1176.150 351.860 ;
        RECT 1175.830 289.920 1176.150 289.980 ;
        RECT 1176.290 289.920 1176.610 289.980 ;
        RECT 1175.830 289.780 1176.610 289.920 ;
        RECT 1175.830 289.720 1176.150 289.780 ;
        RECT 1176.290 289.720 1176.610 289.780 ;
        RECT 1175.830 241.980 1176.150 242.040 ;
        RECT 1176.290 241.980 1176.610 242.040 ;
        RECT 1175.830 241.840 1176.610 241.980 ;
        RECT 1175.830 241.780 1176.150 241.840 ;
        RECT 1176.290 241.780 1176.610 241.840 ;
        RECT 1175.830 234.500 1176.150 234.560 ;
        RECT 1175.635 234.360 1176.150 234.500 ;
        RECT 1175.830 234.300 1176.150 234.360 ;
        RECT 1175.830 186.560 1176.150 186.620 ;
        RECT 1175.635 186.420 1176.150 186.560 ;
        RECT 1175.830 186.360 1176.150 186.420 ;
        RECT 1175.830 96.800 1176.150 96.860 ;
        RECT 1176.290 96.800 1176.610 96.860 ;
        RECT 1175.830 96.660 1176.610 96.800 ;
        RECT 1175.830 96.600 1176.150 96.660 ;
        RECT 1176.290 96.600 1176.610 96.660 ;
        RECT 270.090 18.260 270.410 18.320 ;
        RECT 1175.830 18.260 1176.150 18.320 ;
        RECT 270.090 18.120 1176.150 18.260 ;
        RECT 270.090 18.060 270.410 18.120 ;
        RECT 1175.830 18.060 1176.150 18.120 ;
      LAYER via ;
        RECT 1175.860 1586.820 1176.120 1587.080 ;
        RECT 1176.780 1509.640 1177.040 1509.900 ;
        RECT 1176.780 1490.260 1177.040 1490.520 ;
        RECT 1176.780 1448.780 1177.040 1449.040 ;
        RECT 1175.860 1393.700 1176.120 1393.960 ;
        RECT 1176.780 1393.700 1177.040 1393.960 ;
        RECT 1176.320 1369.560 1176.580 1369.820 ;
        RECT 1175.860 1304.280 1176.120 1304.540 ;
        RECT 1175.860 1296.800 1176.120 1297.060 ;
        RECT 1175.860 1219.960 1176.120 1220.220 ;
        RECT 1174.940 1159.100 1175.200 1159.360 ;
        RECT 1176.320 1159.100 1176.580 1159.360 ;
        RECT 1175.860 1110.820 1176.120 1111.080 ;
        RECT 1176.780 1110.820 1177.040 1111.080 ;
        RECT 1175.860 1013.920 1176.120 1014.180 ;
        RECT 1176.320 1013.920 1176.580 1014.180 ;
        RECT 1176.320 1007.120 1176.580 1007.380 ;
        RECT 1174.940 1006.780 1175.200 1007.040 ;
        RECT 1174.940 917.700 1175.200 917.960 ;
        RECT 1175.860 917.700 1176.120 917.960 ;
        RECT 1174.940 869.420 1175.200 869.680 ;
        RECT 1176.320 869.420 1176.580 869.680 ;
        RECT 1174.940 862.280 1175.200 862.540 ;
        RECT 1176.320 862.280 1176.580 862.540 ;
        RECT 1175.860 813.660 1176.120 813.920 ;
        RECT 1175.860 786.800 1176.120 787.060 ;
        RECT 1175.860 724.240 1176.120 724.500 ;
        RECT 1176.320 723.900 1176.580 724.160 ;
        RECT 1176.320 717.440 1176.580 717.700 ;
        RECT 1176.320 669.500 1176.580 669.760 ;
        RECT 1176.320 620.880 1176.580 621.140 ;
        RECT 1176.320 614.080 1176.580 614.340 ;
        RECT 1176.320 572.260 1176.580 572.520 ;
        RECT 1176.780 572.260 1177.040 572.520 ;
        RECT 1176.780 497.460 1177.040 497.720 ;
        RECT 1175.860 496.780 1176.120 497.040 ;
        RECT 1175.860 434.560 1176.120 434.820 ;
        RECT 1176.320 434.560 1176.580 434.820 ;
        RECT 1176.320 427.420 1176.580 427.680 ;
        RECT 1176.320 379.480 1176.580 379.740 ;
        RECT 1176.320 352.280 1176.580 352.540 ;
        RECT 1175.860 351.600 1176.120 351.860 ;
        RECT 1175.860 289.720 1176.120 289.980 ;
        RECT 1176.320 289.720 1176.580 289.980 ;
        RECT 1175.860 241.780 1176.120 242.040 ;
        RECT 1176.320 241.780 1176.580 242.040 ;
        RECT 1175.860 234.300 1176.120 234.560 ;
        RECT 1175.860 186.360 1176.120 186.620 ;
        RECT 1175.860 96.600 1176.120 96.860 ;
        RECT 1176.320 96.600 1176.580 96.860 ;
        RECT 270.120 18.060 270.380 18.320 ;
        RECT 1175.860 18.060 1176.120 18.320 ;
      LAYER met2 ;
        RECT 1177.140 1700.340 1177.420 1704.000 ;
        RECT 1177.140 1700.000 1177.440 1700.340 ;
        RECT 1177.300 1637.850 1177.440 1700.000 ;
        RECT 1175.920 1637.710 1177.440 1637.850 ;
        RECT 1175.920 1587.110 1176.060 1637.710 ;
        RECT 1175.860 1586.790 1176.120 1587.110 ;
        RECT 1176.780 1509.610 1177.040 1509.930 ;
        RECT 1176.840 1490.550 1176.980 1509.610 ;
        RECT 1176.780 1490.230 1177.040 1490.550 ;
        RECT 1176.780 1448.750 1177.040 1449.070 ;
        RECT 1175.920 1393.990 1176.060 1394.145 ;
        RECT 1176.840 1393.990 1176.980 1448.750 ;
        RECT 1175.860 1393.730 1176.120 1393.990 ;
        RECT 1175.860 1393.670 1176.520 1393.730 ;
        RECT 1176.780 1393.670 1177.040 1393.990 ;
        RECT 1175.920 1393.590 1176.520 1393.670 ;
        RECT 1176.380 1369.850 1176.520 1393.590 ;
        RECT 1176.320 1369.530 1176.580 1369.850 ;
        RECT 1175.860 1304.250 1176.120 1304.570 ;
        RECT 1175.920 1297.090 1176.060 1304.250 ;
        RECT 1175.860 1296.770 1176.120 1297.090 ;
        RECT 1175.860 1219.930 1176.120 1220.250 ;
        RECT 1175.920 1207.525 1176.060 1219.930 ;
        RECT 1174.930 1207.155 1175.210 1207.525 ;
        RECT 1175.850 1207.155 1176.130 1207.525 ;
        RECT 1175.000 1159.390 1175.140 1207.155 ;
        RECT 1174.940 1159.070 1175.200 1159.390 ;
        RECT 1176.320 1159.070 1176.580 1159.390 ;
        RECT 1176.380 1125.130 1176.520 1159.070 ;
        RECT 1176.380 1124.990 1176.980 1125.130 ;
        RECT 1176.840 1111.110 1176.980 1124.990 ;
        RECT 1175.860 1110.790 1176.120 1111.110 ;
        RECT 1176.780 1110.790 1177.040 1111.110 ;
        RECT 1175.920 1104.165 1176.060 1110.790 ;
        RECT 1174.930 1103.795 1175.210 1104.165 ;
        RECT 1175.850 1103.795 1176.130 1104.165 ;
        RECT 1175.000 1055.885 1175.140 1103.795 ;
        RECT 1174.930 1055.515 1175.210 1055.885 ;
        RECT 1175.850 1055.515 1176.130 1055.885 ;
        RECT 1175.920 1014.210 1176.060 1055.515 ;
        RECT 1175.860 1013.890 1176.120 1014.210 ;
        RECT 1176.320 1013.890 1176.580 1014.210 ;
        RECT 1176.380 1007.410 1176.520 1013.890 ;
        RECT 1176.320 1007.090 1176.580 1007.410 ;
        RECT 1174.940 1006.750 1175.200 1007.070 ;
        RECT 1175.000 917.990 1175.140 1006.750 ;
        RECT 1174.940 917.845 1175.200 917.990 ;
        RECT 1175.860 917.845 1176.120 917.990 ;
        RECT 1174.930 917.475 1175.210 917.845 ;
        RECT 1175.850 917.475 1176.130 917.845 ;
        RECT 1175.000 869.710 1175.140 917.475 ;
        RECT 1174.940 869.390 1175.200 869.710 ;
        RECT 1176.320 869.390 1176.580 869.710 ;
        RECT 1176.380 862.570 1176.520 869.390 ;
        RECT 1174.940 862.250 1175.200 862.570 ;
        RECT 1176.320 862.250 1176.580 862.570 ;
        RECT 1175.000 814.485 1175.140 862.250 ;
        RECT 1174.930 814.115 1175.210 814.485 ;
        RECT 1175.850 814.115 1176.130 814.485 ;
        RECT 1175.920 813.950 1176.060 814.115 ;
        RECT 1175.860 813.630 1176.120 813.950 ;
        RECT 1175.860 786.770 1176.120 787.090 ;
        RECT 1175.920 724.530 1176.060 786.770 ;
        RECT 1175.860 724.210 1176.120 724.530 ;
        RECT 1176.320 723.870 1176.580 724.190 ;
        RECT 1176.380 717.730 1176.520 723.870 ;
        RECT 1176.320 717.410 1176.580 717.730 ;
        RECT 1176.320 669.470 1176.580 669.790 ;
        RECT 1176.380 621.170 1176.520 669.470 ;
        RECT 1176.320 620.850 1176.580 621.170 ;
        RECT 1176.320 614.050 1176.580 614.370 ;
        RECT 1176.380 572.550 1176.520 614.050 ;
        RECT 1176.320 572.230 1176.580 572.550 ;
        RECT 1176.780 572.230 1177.040 572.550 ;
        RECT 1176.840 497.750 1176.980 572.230 ;
        RECT 1176.780 497.430 1177.040 497.750 ;
        RECT 1175.860 496.750 1176.120 497.070 ;
        RECT 1175.920 434.850 1176.060 496.750 ;
        RECT 1175.860 434.530 1176.120 434.850 ;
        RECT 1176.320 434.530 1176.580 434.850 ;
        RECT 1176.380 427.710 1176.520 434.530 ;
        RECT 1176.320 427.390 1176.580 427.710 ;
        RECT 1176.320 379.450 1176.580 379.770 ;
        RECT 1176.380 352.570 1176.520 379.450 ;
        RECT 1176.320 352.250 1176.580 352.570 ;
        RECT 1175.860 351.570 1176.120 351.890 ;
        RECT 1175.920 290.010 1176.060 351.570 ;
        RECT 1175.860 289.690 1176.120 290.010 ;
        RECT 1176.320 289.690 1176.580 290.010 ;
        RECT 1176.380 242.070 1176.520 289.690 ;
        RECT 1175.860 241.750 1176.120 242.070 ;
        RECT 1176.320 241.750 1176.580 242.070 ;
        RECT 1175.920 234.590 1176.060 241.750 ;
        RECT 1175.860 234.270 1176.120 234.590 ;
        RECT 1175.860 186.330 1176.120 186.650 ;
        RECT 1175.920 96.890 1176.060 186.330 ;
        RECT 1175.860 96.570 1176.120 96.890 ;
        RECT 1176.320 96.570 1176.580 96.890 ;
        RECT 1176.380 72.490 1176.520 96.570 ;
        RECT 1175.920 72.350 1176.520 72.490 ;
        RECT 1175.920 18.350 1176.060 72.350 ;
        RECT 270.120 18.030 270.380 18.350 ;
        RECT 1175.860 18.030 1176.120 18.350 ;
        RECT 270.180 2.400 270.320 18.030 ;
        RECT 269.970 -4.800 270.530 2.400 ;
      LAYER via2 ;
        RECT 1174.930 1207.200 1175.210 1207.480 ;
        RECT 1175.850 1207.200 1176.130 1207.480 ;
        RECT 1174.930 1103.840 1175.210 1104.120 ;
        RECT 1175.850 1103.840 1176.130 1104.120 ;
        RECT 1174.930 1055.560 1175.210 1055.840 ;
        RECT 1175.850 1055.560 1176.130 1055.840 ;
        RECT 1174.930 917.520 1175.210 917.800 ;
        RECT 1175.850 917.520 1176.130 917.800 ;
        RECT 1174.930 814.160 1175.210 814.440 ;
        RECT 1175.850 814.160 1176.130 814.440 ;
      LAYER met3 ;
        RECT 1174.905 1207.490 1175.235 1207.505 ;
        RECT 1175.825 1207.490 1176.155 1207.505 ;
        RECT 1174.905 1207.190 1176.155 1207.490 ;
        RECT 1174.905 1207.175 1175.235 1207.190 ;
        RECT 1175.825 1207.175 1176.155 1207.190 ;
        RECT 1174.905 1104.130 1175.235 1104.145 ;
        RECT 1175.825 1104.130 1176.155 1104.145 ;
        RECT 1174.905 1103.830 1176.155 1104.130 ;
        RECT 1174.905 1103.815 1175.235 1103.830 ;
        RECT 1175.825 1103.815 1176.155 1103.830 ;
        RECT 1174.905 1055.850 1175.235 1055.865 ;
        RECT 1175.825 1055.850 1176.155 1055.865 ;
        RECT 1174.905 1055.550 1176.155 1055.850 ;
        RECT 1174.905 1055.535 1175.235 1055.550 ;
        RECT 1175.825 1055.535 1176.155 1055.550 ;
        RECT 1174.905 917.810 1175.235 917.825 ;
        RECT 1175.825 917.810 1176.155 917.825 ;
        RECT 1174.905 917.510 1176.155 917.810 ;
        RECT 1174.905 917.495 1175.235 917.510 ;
        RECT 1175.825 917.495 1176.155 917.510 ;
        RECT 1174.905 814.450 1175.235 814.465 ;
        RECT 1175.825 814.450 1176.155 814.465 ;
        RECT 1174.905 814.150 1176.155 814.450 ;
        RECT 1174.905 814.135 1175.235 814.150 ;
        RECT 1175.825 814.135 1176.155 814.150 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1177.745 1352.605 1177.915 1400.715 ;
        RECT 1177.745 676.345 1177.915 724.455 ;
        RECT 1177.745 579.785 1177.915 627.895 ;
        RECT 1177.745 289.765 1177.915 337.875 ;
        RECT 1177.745 96.645 1177.915 144.755 ;
        RECT 1148.765 18.445 1148.935 19.295 ;
      LAYER mcon ;
        RECT 1177.745 1400.545 1177.915 1400.715 ;
        RECT 1177.745 724.285 1177.915 724.455 ;
        RECT 1177.745 627.725 1177.915 627.895 ;
        RECT 1177.745 337.705 1177.915 337.875 ;
        RECT 1177.745 144.585 1177.915 144.755 ;
        RECT 1148.765 19.125 1148.935 19.295 ;
      LAYER met1 ;
        RECT 1177.670 1658.080 1177.990 1658.140 ;
        RECT 1179.050 1658.080 1179.370 1658.140 ;
        RECT 1177.670 1657.940 1179.370 1658.080 ;
        RECT 1177.670 1657.880 1177.990 1657.940 ;
        RECT 1179.050 1657.880 1179.370 1657.940 ;
        RECT 1177.670 1400.700 1177.990 1400.760 ;
        RECT 1177.475 1400.560 1177.990 1400.700 ;
        RECT 1177.670 1400.500 1177.990 1400.560 ;
        RECT 1177.670 1352.760 1177.990 1352.820 ;
        RECT 1177.475 1352.620 1177.990 1352.760 ;
        RECT 1177.670 1352.560 1177.990 1352.620 ;
        RECT 1177.670 1152.500 1177.990 1152.560 ;
        RECT 1178.590 1152.500 1178.910 1152.560 ;
        RECT 1177.670 1152.360 1178.910 1152.500 ;
        RECT 1177.670 1152.300 1177.990 1152.360 ;
        RECT 1178.590 1152.300 1178.910 1152.360 ;
        RECT 1177.670 1014.460 1177.990 1014.520 ;
        RECT 1178.130 1014.460 1178.450 1014.520 ;
        RECT 1177.670 1014.320 1178.450 1014.460 ;
        RECT 1177.670 1014.260 1177.990 1014.320 ;
        RECT 1178.130 1014.260 1178.450 1014.320 ;
        RECT 1177.670 966.180 1177.990 966.240 ;
        RECT 1178.130 966.180 1178.450 966.240 ;
        RECT 1177.670 966.040 1178.450 966.180 ;
        RECT 1177.670 965.980 1177.990 966.040 ;
        RECT 1178.130 965.980 1178.450 966.040 ;
        RECT 1177.210 869.620 1177.530 869.680 ;
        RECT 1177.670 869.620 1177.990 869.680 ;
        RECT 1177.210 869.480 1177.990 869.620 ;
        RECT 1177.210 869.420 1177.530 869.480 ;
        RECT 1177.670 869.420 1177.990 869.480 ;
        RECT 1177.670 724.440 1177.990 724.500 ;
        RECT 1177.475 724.300 1177.990 724.440 ;
        RECT 1177.670 724.240 1177.990 724.300 ;
        RECT 1177.670 676.500 1177.990 676.560 ;
        RECT 1177.475 676.360 1177.990 676.500 ;
        RECT 1177.670 676.300 1177.990 676.360 ;
        RECT 1177.670 627.880 1177.990 627.940 ;
        RECT 1177.475 627.740 1177.990 627.880 ;
        RECT 1177.670 627.680 1177.990 627.740 ;
        RECT 1177.670 579.940 1177.990 580.000 ;
        RECT 1177.475 579.800 1177.990 579.940 ;
        RECT 1177.670 579.740 1177.990 579.800 ;
        RECT 1177.210 386.480 1177.530 386.540 ;
        RECT 1177.670 386.480 1177.990 386.540 ;
        RECT 1177.210 386.340 1177.990 386.480 ;
        RECT 1177.210 386.280 1177.530 386.340 ;
        RECT 1177.670 386.280 1177.990 386.340 ;
        RECT 1177.670 337.860 1177.990 337.920 ;
        RECT 1177.475 337.720 1177.990 337.860 ;
        RECT 1177.670 337.660 1177.990 337.720 ;
        RECT 1177.670 289.920 1177.990 289.980 ;
        RECT 1177.475 289.780 1177.990 289.920 ;
        RECT 1177.670 289.720 1177.990 289.780 ;
        RECT 1177.670 144.740 1177.990 144.800 ;
        RECT 1177.475 144.600 1177.990 144.740 ;
        RECT 1177.670 144.540 1177.990 144.600 ;
        RECT 1177.670 96.800 1177.990 96.860 ;
        RECT 1177.475 96.660 1177.990 96.800 ;
        RECT 1177.670 96.600 1177.990 96.660 ;
        RECT 1148.705 19.280 1148.995 19.325 ;
        RECT 1177.670 19.280 1177.990 19.340 ;
        RECT 1148.705 19.140 1177.990 19.280 ;
        RECT 1148.705 19.095 1148.995 19.140 ;
        RECT 1177.670 19.080 1177.990 19.140 ;
        RECT 288.030 18.600 288.350 18.660 ;
        RECT 1148.705 18.600 1148.995 18.645 ;
        RECT 288.030 18.460 1148.995 18.600 ;
        RECT 288.030 18.400 288.350 18.460 ;
        RECT 1148.705 18.415 1148.995 18.460 ;
      LAYER via ;
        RECT 1177.700 1657.880 1177.960 1658.140 ;
        RECT 1179.080 1657.880 1179.340 1658.140 ;
        RECT 1177.700 1400.500 1177.960 1400.760 ;
        RECT 1177.700 1352.560 1177.960 1352.820 ;
        RECT 1177.700 1152.300 1177.960 1152.560 ;
        RECT 1178.620 1152.300 1178.880 1152.560 ;
        RECT 1177.700 1014.260 1177.960 1014.520 ;
        RECT 1178.160 1014.260 1178.420 1014.520 ;
        RECT 1177.700 965.980 1177.960 966.240 ;
        RECT 1178.160 965.980 1178.420 966.240 ;
        RECT 1177.240 869.420 1177.500 869.680 ;
        RECT 1177.700 869.420 1177.960 869.680 ;
        RECT 1177.700 724.240 1177.960 724.500 ;
        RECT 1177.700 676.300 1177.960 676.560 ;
        RECT 1177.700 627.680 1177.960 627.940 ;
        RECT 1177.700 579.740 1177.960 580.000 ;
        RECT 1177.240 386.280 1177.500 386.540 ;
        RECT 1177.700 386.280 1177.960 386.540 ;
        RECT 1177.700 337.660 1177.960 337.920 ;
        RECT 1177.700 289.720 1177.960 289.980 ;
        RECT 1177.700 144.540 1177.960 144.800 ;
        RECT 1177.700 96.600 1177.960 96.860 ;
        RECT 1177.700 19.080 1177.960 19.340 ;
        RECT 288.060 18.400 288.320 18.660 ;
      LAYER met2 ;
        RECT 1178.980 1700.340 1179.260 1704.000 ;
        RECT 1178.980 1700.000 1179.280 1700.340 ;
        RECT 1179.140 1658.170 1179.280 1700.000 ;
        RECT 1177.700 1657.850 1177.960 1658.170 ;
        RECT 1179.080 1657.850 1179.340 1658.170 ;
        RECT 1177.760 1400.790 1177.900 1657.850 ;
        RECT 1177.700 1400.470 1177.960 1400.790 ;
        RECT 1177.700 1352.530 1177.960 1352.850 ;
        RECT 1177.760 1207.525 1177.900 1352.530 ;
        RECT 1177.690 1207.155 1177.970 1207.525 ;
        RECT 1178.610 1207.155 1178.890 1207.525 ;
        RECT 1178.680 1152.590 1178.820 1207.155 ;
        RECT 1177.700 1152.270 1177.960 1152.590 ;
        RECT 1178.620 1152.270 1178.880 1152.590 ;
        RECT 1177.760 1104.165 1177.900 1152.270 ;
        RECT 1177.690 1103.795 1177.970 1104.165 ;
        RECT 1178.610 1103.795 1178.890 1104.165 ;
        RECT 1178.680 1055.885 1178.820 1103.795 ;
        RECT 1177.690 1055.515 1177.970 1055.885 ;
        RECT 1178.610 1055.515 1178.890 1055.885 ;
        RECT 1177.760 1014.550 1177.900 1055.515 ;
        RECT 1177.700 1014.230 1177.960 1014.550 ;
        RECT 1178.160 1014.230 1178.420 1014.550 ;
        RECT 1178.220 966.270 1178.360 1014.230 ;
        RECT 1177.700 965.950 1177.960 966.270 ;
        RECT 1178.160 965.950 1178.420 966.270 ;
        RECT 1177.760 942.210 1177.900 965.950 ;
        RECT 1177.300 942.070 1177.900 942.210 ;
        RECT 1177.300 869.710 1177.440 942.070 ;
        RECT 1177.240 869.390 1177.500 869.710 ;
        RECT 1177.700 869.390 1177.960 869.710 ;
        RECT 1177.760 724.530 1177.900 869.390 ;
        RECT 1177.700 724.210 1177.960 724.530 ;
        RECT 1177.700 676.270 1177.960 676.590 ;
        RECT 1177.760 627.970 1177.900 676.270 ;
        RECT 1177.700 627.650 1177.960 627.970 ;
        RECT 1177.700 579.710 1177.960 580.030 ;
        RECT 1177.760 435.725 1177.900 579.710 ;
        RECT 1177.690 435.355 1177.970 435.725 ;
        RECT 1177.230 434.675 1177.510 435.045 ;
        RECT 1177.300 386.570 1177.440 434.675 ;
        RECT 1177.240 386.250 1177.500 386.570 ;
        RECT 1177.700 386.250 1177.960 386.570 ;
        RECT 1177.760 337.950 1177.900 386.250 ;
        RECT 1177.700 337.630 1177.960 337.950 ;
        RECT 1177.700 289.690 1177.960 290.010 ;
        RECT 1177.760 144.830 1177.900 289.690 ;
        RECT 1177.700 144.510 1177.960 144.830 ;
        RECT 1177.700 96.570 1177.960 96.890 ;
        RECT 1177.760 19.370 1177.900 96.570 ;
        RECT 1177.700 19.050 1177.960 19.370 ;
        RECT 288.060 18.370 288.320 18.690 ;
        RECT 288.120 2.400 288.260 18.370 ;
        RECT 287.910 -4.800 288.470 2.400 ;
      LAYER via2 ;
        RECT 1177.690 1207.200 1177.970 1207.480 ;
        RECT 1178.610 1207.200 1178.890 1207.480 ;
        RECT 1177.690 1103.840 1177.970 1104.120 ;
        RECT 1178.610 1103.840 1178.890 1104.120 ;
        RECT 1177.690 1055.560 1177.970 1055.840 ;
        RECT 1178.610 1055.560 1178.890 1055.840 ;
        RECT 1177.690 435.400 1177.970 435.680 ;
        RECT 1177.230 434.720 1177.510 435.000 ;
      LAYER met3 ;
        RECT 1177.665 1207.490 1177.995 1207.505 ;
        RECT 1178.585 1207.490 1178.915 1207.505 ;
        RECT 1177.665 1207.190 1178.915 1207.490 ;
        RECT 1177.665 1207.175 1177.995 1207.190 ;
        RECT 1178.585 1207.175 1178.915 1207.190 ;
        RECT 1177.665 1104.130 1177.995 1104.145 ;
        RECT 1178.585 1104.130 1178.915 1104.145 ;
        RECT 1177.665 1103.830 1178.915 1104.130 ;
        RECT 1177.665 1103.815 1177.995 1103.830 ;
        RECT 1178.585 1103.815 1178.915 1103.830 ;
        RECT 1177.665 1055.850 1177.995 1055.865 ;
        RECT 1178.585 1055.850 1178.915 1055.865 ;
        RECT 1177.665 1055.550 1178.915 1055.850 ;
        RECT 1177.665 1055.535 1177.995 1055.550 ;
        RECT 1178.585 1055.535 1178.915 1055.550 ;
        RECT 1177.665 435.690 1177.995 435.705 ;
        RECT 1176.990 435.390 1177.995 435.690 ;
        RECT 1176.990 435.025 1177.290 435.390 ;
        RECT 1177.665 435.375 1177.995 435.390 ;
        RECT 1176.990 434.710 1177.535 435.025 ;
        RECT 1177.205 434.695 1177.535 434.710 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 305.970 18.940 306.290 19.000 ;
        RECT 1180.430 18.940 1180.750 19.000 ;
        RECT 305.970 18.800 1180.750 18.940 ;
        RECT 305.970 18.740 306.290 18.800 ;
        RECT 1180.430 18.740 1180.750 18.800 ;
      LAYER via ;
        RECT 306.000 18.740 306.260 19.000 ;
        RECT 1180.460 18.740 1180.720 19.000 ;
      LAYER met2 ;
        RECT 1180.820 1700.340 1181.100 1704.000 ;
        RECT 1180.820 1700.000 1181.120 1700.340 ;
        RECT 1180.980 1677.290 1181.120 1700.000 ;
        RECT 1180.520 1677.150 1181.120 1677.290 ;
        RECT 1180.520 19.030 1180.660 1677.150 ;
        RECT 306.000 18.710 306.260 19.030 ;
        RECT 1180.460 18.710 1180.720 19.030 ;
        RECT 306.060 2.400 306.200 18.710 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1185.105 1594.005 1185.275 1642.115 ;
        RECT 1186.025 1490.645 1186.195 1538.755 ;
        RECT 1185.565 1207.425 1185.735 1255.875 ;
        RECT 1185.105 379.865 1185.275 427.635 ;
        RECT 1186.025 289.765 1186.195 379.355 ;
        RECT 1126.225 17.425 1126.395 19.295 ;
        RECT 1148.305 16.745 1148.475 17.595 ;
      LAYER mcon ;
        RECT 1185.105 1641.945 1185.275 1642.115 ;
        RECT 1186.025 1538.585 1186.195 1538.755 ;
        RECT 1185.565 1255.705 1185.735 1255.875 ;
        RECT 1185.105 427.465 1185.275 427.635 ;
        RECT 1186.025 379.185 1186.195 379.355 ;
        RECT 1126.225 19.125 1126.395 19.295 ;
        RECT 1148.305 17.425 1148.475 17.595 ;
      LAYER met1 ;
        RECT 1182.730 1680.520 1183.050 1680.580 ;
        RECT 1184.570 1680.520 1184.890 1680.580 ;
        RECT 1182.730 1680.380 1184.890 1680.520 ;
        RECT 1182.730 1680.320 1183.050 1680.380 ;
        RECT 1184.570 1680.320 1184.890 1680.380 ;
        RECT 1185.030 1642.100 1185.350 1642.160 ;
        RECT 1184.835 1641.960 1185.350 1642.100 ;
        RECT 1185.030 1641.900 1185.350 1641.960 ;
        RECT 1185.045 1594.160 1185.335 1594.205 ;
        RECT 1185.490 1594.160 1185.810 1594.220 ;
        RECT 1185.045 1594.020 1185.810 1594.160 ;
        RECT 1185.045 1593.975 1185.335 1594.020 ;
        RECT 1185.490 1593.960 1185.810 1594.020 ;
        RECT 1185.965 1538.740 1186.255 1538.785 ;
        RECT 1186.410 1538.740 1186.730 1538.800 ;
        RECT 1185.965 1538.600 1186.730 1538.740 ;
        RECT 1185.965 1538.555 1186.255 1538.600 ;
        RECT 1186.410 1538.540 1186.730 1538.600 ;
        RECT 1185.950 1490.800 1186.270 1490.860 ;
        RECT 1185.755 1490.660 1186.270 1490.800 ;
        RECT 1185.950 1490.600 1186.270 1490.660 ;
        RECT 1185.490 1400.700 1185.810 1400.760 ;
        RECT 1185.950 1400.700 1186.270 1400.760 ;
        RECT 1185.490 1400.560 1186.270 1400.700 ;
        RECT 1185.490 1400.500 1185.810 1400.560 ;
        RECT 1185.950 1400.500 1186.270 1400.560 ;
        RECT 1185.030 1269.460 1185.350 1269.520 ;
        RECT 1185.950 1269.460 1186.270 1269.520 ;
        RECT 1185.030 1269.320 1186.270 1269.460 ;
        RECT 1185.030 1269.260 1185.350 1269.320 ;
        RECT 1185.950 1269.260 1186.270 1269.320 ;
        RECT 1185.505 1255.860 1185.795 1255.905 ;
        RECT 1185.950 1255.860 1186.270 1255.920 ;
        RECT 1185.505 1255.720 1186.270 1255.860 ;
        RECT 1185.505 1255.675 1185.795 1255.720 ;
        RECT 1185.950 1255.660 1186.270 1255.720 ;
        RECT 1185.490 1207.580 1185.810 1207.640 ;
        RECT 1185.295 1207.440 1185.810 1207.580 ;
        RECT 1185.490 1207.380 1185.810 1207.440 ;
        RECT 1185.030 1062.540 1185.350 1062.800 ;
        RECT 1185.120 1062.120 1185.260 1062.540 ;
        RECT 1185.030 1061.860 1185.350 1062.120 ;
        RECT 1185.490 1014.120 1185.810 1014.180 ;
        RECT 1185.950 1014.120 1186.270 1014.180 ;
        RECT 1185.490 1013.980 1186.270 1014.120 ;
        RECT 1185.490 1013.920 1185.810 1013.980 ;
        RECT 1185.950 1013.920 1186.270 1013.980 ;
        RECT 1185.490 917.560 1185.810 917.620 ;
        RECT 1185.950 917.560 1186.270 917.620 ;
        RECT 1185.490 917.420 1186.270 917.560 ;
        RECT 1185.490 917.360 1185.810 917.420 ;
        RECT 1185.950 917.360 1186.270 917.420 ;
        RECT 1185.030 786.660 1185.350 786.720 ;
        RECT 1185.950 786.660 1186.270 786.720 ;
        RECT 1185.030 786.520 1186.270 786.660 ;
        RECT 1185.030 786.460 1185.350 786.520 ;
        RECT 1185.950 786.460 1186.270 786.520 ;
        RECT 1185.490 724.780 1185.810 724.840 ;
        RECT 1185.950 724.780 1186.270 724.840 ;
        RECT 1185.490 724.640 1186.270 724.780 ;
        RECT 1185.490 724.580 1185.810 724.640 ;
        RECT 1185.950 724.580 1186.270 724.640 ;
        RECT 1185.490 689.900 1185.810 690.160 ;
        RECT 1185.580 689.760 1185.720 689.900 ;
        RECT 1185.950 689.760 1186.270 689.820 ;
        RECT 1185.580 689.620 1186.270 689.760 ;
        RECT 1185.950 689.560 1186.270 689.620 ;
        RECT 1185.490 593.340 1185.810 593.600 ;
        RECT 1185.580 593.200 1185.720 593.340 ;
        RECT 1185.950 593.200 1186.270 593.260 ;
        RECT 1185.580 593.060 1186.270 593.200 ;
        RECT 1185.950 593.000 1186.270 593.060 ;
        RECT 1185.045 427.620 1185.335 427.665 ;
        RECT 1185.950 427.620 1186.270 427.680 ;
        RECT 1185.045 427.480 1186.270 427.620 ;
        RECT 1185.045 427.435 1185.335 427.480 ;
        RECT 1185.950 427.420 1186.270 427.480 ;
        RECT 1185.030 380.020 1185.350 380.080 ;
        RECT 1184.835 379.880 1185.350 380.020 ;
        RECT 1185.030 379.820 1185.350 379.880 ;
        RECT 1185.030 379.340 1185.350 379.400 ;
        RECT 1185.965 379.340 1186.255 379.385 ;
        RECT 1185.030 379.200 1186.255 379.340 ;
        RECT 1185.030 379.140 1185.350 379.200 ;
        RECT 1185.965 379.155 1186.255 379.200 ;
        RECT 1185.950 289.920 1186.270 289.980 ;
        RECT 1185.755 289.780 1186.270 289.920 ;
        RECT 1185.950 289.720 1186.270 289.780 ;
        RECT 1185.950 255.580 1186.270 255.640 ;
        RECT 1185.580 255.440 1186.270 255.580 ;
        RECT 1185.580 255.300 1185.720 255.440 ;
        RECT 1185.950 255.380 1186.270 255.440 ;
        RECT 1185.490 255.040 1185.810 255.300 ;
        RECT 1185.030 206.960 1185.350 207.020 ;
        RECT 1185.950 206.960 1186.270 207.020 ;
        RECT 1185.030 206.820 1186.270 206.960 ;
        RECT 1185.030 206.760 1185.350 206.820 ;
        RECT 1185.950 206.760 1186.270 206.820 ;
        RECT 1185.950 159.020 1186.270 159.080 ;
        RECT 1185.120 158.880 1186.270 159.020 ;
        RECT 1185.120 158.740 1185.260 158.880 ;
        RECT 1185.950 158.820 1186.270 158.880 ;
        RECT 1185.030 158.480 1185.350 158.740 ;
        RECT 1185.030 96.800 1185.350 96.860 ;
        RECT 1185.490 96.800 1185.810 96.860 ;
        RECT 1185.030 96.660 1185.810 96.800 ;
        RECT 1185.030 96.600 1185.350 96.660 ;
        RECT 1185.490 96.600 1185.810 96.660 ;
        RECT 323.450 19.280 323.770 19.340 ;
        RECT 1126.165 19.280 1126.455 19.325 ;
        RECT 323.450 19.140 1126.455 19.280 ;
        RECT 323.450 19.080 323.770 19.140 ;
        RECT 1126.165 19.095 1126.455 19.140 ;
        RECT 1126.165 17.580 1126.455 17.625 ;
        RECT 1148.245 17.580 1148.535 17.625 ;
        RECT 1126.165 17.440 1148.535 17.580 ;
        RECT 1126.165 17.395 1126.455 17.440 ;
        RECT 1148.245 17.395 1148.535 17.440 ;
        RECT 1148.245 16.900 1148.535 16.945 ;
        RECT 1185.030 16.900 1185.350 16.960 ;
        RECT 1148.245 16.760 1185.350 16.900 ;
        RECT 1148.245 16.715 1148.535 16.760 ;
        RECT 1185.030 16.700 1185.350 16.760 ;
      LAYER via ;
        RECT 1182.760 1680.320 1183.020 1680.580 ;
        RECT 1184.600 1680.320 1184.860 1680.580 ;
        RECT 1185.060 1641.900 1185.320 1642.160 ;
        RECT 1185.520 1593.960 1185.780 1594.220 ;
        RECT 1186.440 1538.540 1186.700 1538.800 ;
        RECT 1185.980 1490.600 1186.240 1490.860 ;
        RECT 1185.520 1400.500 1185.780 1400.760 ;
        RECT 1185.980 1400.500 1186.240 1400.760 ;
        RECT 1185.060 1269.260 1185.320 1269.520 ;
        RECT 1185.980 1269.260 1186.240 1269.520 ;
        RECT 1185.980 1255.660 1186.240 1255.920 ;
        RECT 1185.520 1207.380 1185.780 1207.640 ;
        RECT 1185.060 1062.540 1185.320 1062.800 ;
        RECT 1185.060 1061.860 1185.320 1062.120 ;
        RECT 1185.520 1013.920 1185.780 1014.180 ;
        RECT 1185.980 1013.920 1186.240 1014.180 ;
        RECT 1185.520 917.360 1185.780 917.620 ;
        RECT 1185.980 917.360 1186.240 917.620 ;
        RECT 1185.060 786.460 1185.320 786.720 ;
        RECT 1185.980 786.460 1186.240 786.720 ;
        RECT 1185.520 724.580 1185.780 724.840 ;
        RECT 1185.980 724.580 1186.240 724.840 ;
        RECT 1185.520 689.900 1185.780 690.160 ;
        RECT 1185.980 689.560 1186.240 689.820 ;
        RECT 1185.520 593.340 1185.780 593.600 ;
        RECT 1185.980 593.000 1186.240 593.260 ;
        RECT 1185.980 427.420 1186.240 427.680 ;
        RECT 1185.060 379.820 1185.320 380.080 ;
        RECT 1185.060 379.140 1185.320 379.400 ;
        RECT 1185.980 289.720 1186.240 289.980 ;
        RECT 1185.980 255.380 1186.240 255.640 ;
        RECT 1185.520 255.040 1185.780 255.300 ;
        RECT 1185.060 206.760 1185.320 207.020 ;
        RECT 1185.980 206.760 1186.240 207.020 ;
        RECT 1185.980 158.820 1186.240 159.080 ;
        RECT 1185.060 158.480 1185.320 158.740 ;
        RECT 1185.060 96.600 1185.320 96.860 ;
        RECT 1185.520 96.600 1185.780 96.860 ;
        RECT 323.480 19.080 323.740 19.340 ;
        RECT 1185.060 16.700 1185.320 16.960 ;
      LAYER met2 ;
        RECT 1182.660 1700.340 1182.940 1704.000 ;
        RECT 1182.660 1700.000 1182.960 1700.340 ;
        RECT 1182.820 1680.610 1182.960 1700.000 ;
        RECT 1182.760 1680.290 1183.020 1680.610 ;
        RECT 1184.600 1680.290 1184.860 1680.610 ;
        RECT 1184.660 1677.460 1184.800 1680.290 ;
        RECT 1184.660 1677.320 1185.260 1677.460 ;
        RECT 1185.120 1642.190 1185.260 1677.320 ;
        RECT 1185.060 1641.870 1185.320 1642.190 ;
        RECT 1185.520 1593.930 1185.780 1594.250 ;
        RECT 1185.580 1562.880 1185.720 1593.930 ;
        RECT 1185.580 1562.740 1186.640 1562.880 ;
        RECT 1186.500 1538.830 1186.640 1562.740 ;
        RECT 1186.440 1538.510 1186.700 1538.830 ;
        RECT 1185.980 1490.570 1186.240 1490.890 ;
        RECT 1186.040 1414.130 1186.180 1490.570 ;
        RECT 1185.580 1413.990 1186.180 1414.130 ;
        RECT 1185.580 1400.790 1185.720 1413.990 ;
        RECT 1185.520 1400.470 1185.780 1400.790 ;
        RECT 1185.980 1400.470 1186.240 1400.790 ;
        RECT 1186.040 1317.570 1186.180 1400.470 ;
        RECT 1185.580 1317.430 1186.180 1317.570 ;
        RECT 1185.580 1269.970 1185.720 1317.430 ;
        RECT 1185.120 1269.830 1185.720 1269.970 ;
        RECT 1185.120 1269.550 1185.260 1269.830 ;
        RECT 1185.060 1269.230 1185.320 1269.550 ;
        RECT 1185.980 1269.230 1186.240 1269.550 ;
        RECT 1186.040 1255.950 1186.180 1269.230 ;
        RECT 1185.980 1255.630 1186.240 1255.950 ;
        RECT 1185.520 1207.350 1185.780 1207.670 ;
        RECT 1185.580 1104.050 1185.720 1207.350 ;
        RECT 1185.120 1103.910 1185.720 1104.050 ;
        RECT 1185.120 1062.830 1185.260 1103.910 ;
        RECT 1185.060 1062.510 1185.320 1062.830 ;
        RECT 1185.060 1061.830 1185.320 1062.150 ;
        RECT 1185.120 1027.890 1185.260 1061.830 ;
        RECT 1185.120 1027.750 1185.720 1027.890 ;
        RECT 1185.580 1014.210 1185.720 1027.750 ;
        RECT 1185.520 1013.890 1185.780 1014.210 ;
        RECT 1185.980 1013.890 1186.240 1014.210 ;
        RECT 1186.040 931.330 1186.180 1013.890 ;
        RECT 1185.580 931.190 1186.180 931.330 ;
        RECT 1185.580 917.650 1185.720 931.190 ;
        RECT 1185.520 917.330 1185.780 917.650 ;
        RECT 1185.980 917.330 1186.240 917.650 ;
        RECT 1186.040 834.770 1186.180 917.330 ;
        RECT 1185.580 834.630 1186.180 834.770 ;
        RECT 1185.580 787.170 1185.720 834.630 ;
        RECT 1185.120 787.030 1185.720 787.170 ;
        RECT 1185.120 786.750 1185.260 787.030 ;
        RECT 1185.060 786.430 1185.320 786.750 ;
        RECT 1185.980 786.430 1186.240 786.750 ;
        RECT 1186.040 724.870 1186.180 786.430 ;
        RECT 1185.520 724.550 1185.780 724.870 ;
        RECT 1185.980 724.550 1186.240 724.870 ;
        RECT 1185.580 690.190 1185.720 724.550 ;
        RECT 1185.520 689.870 1185.780 690.190 ;
        RECT 1185.980 689.530 1186.240 689.850 ;
        RECT 1186.040 641.650 1186.180 689.530 ;
        RECT 1185.580 641.510 1186.180 641.650 ;
        RECT 1185.580 593.630 1185.720 641.510 ;
        RECT 1185.520 593.310 1185.780 593.630 ;
        RECT 1185.980 592.970 1186.240 593.290 ;
        RECT 1186.040 545.090 1186.180 592.970 ;
        RECT 1185.580 544.950 1186.180 545.090 ;
        RECT 1185.580 500.210 1185.720 544.950 ;
        RECT 1185.580 500.070 1186.180 500.210 ;
        RECT 1186.040 427.710 1186.180 500.070 ;
        RECT 1185.980 427.390 1186.240 427.710 ;
        RECT 1185.060 379.790 1185.320 380.110 ;
        RECT 1185.120 379.430 1185.260 379.790 ;
        RECT 1185.060 379.110 1185.320 379.430 ;
        RECT 1185.980 289.690 1186.240 290.010 ;
        RECT 1186.040 255.670 1186.180 289.690 ;
        RECT 1185.980 255.350 1186.240 255.670 ;
        RECT 1185.520 255.010 1185.780 255.330 ;
        RECT 1185.580 207.130 1185.720 255.010 ;
        RECT 1185.120 207.050 1185.720 207.130 ;
        RECT 1185.060 206.990 1185.720 207.050 ;
        RECT 1185.060 206.730 1185.320 206.990 ;
        RECT 1185.980 206.730 1186.240 207.050 ;
        RECT 1186.040 159.110 1186.180 206.730 ;
        RECT 1185.980 158.790 1186.240 159.110 ;
        RECT 1185.060 158.450 1185.320 158.770 ;
        RECT 1185.120 96.890 1185.260 158.450 ;
        RECT 1185.060 96.570 1185.320 96.890 ;
        RECT 1185.520 96.570 1185.780 96.890 ;
        RECT 1185.580 72.490 1185.720 96.570 ;
        RECT 1185.120 72.350 1185.720 72.490 ;
        RECT 323.480 19.050 323.740 19.370 ;
        RECT 323.540 9.930 323.680 19.050 ;
        RECT 1185.120 16.990 1185.260 72.350 ;
        RECT 1185.060 16.670 1185.320 16.990 ;
        RECT 323.540 9.790 324.140 9.930 ;
        RECT 324.000 2.400 324.140 9.790 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1180.890 1676.780 1181.210 1676.840 ;
        RECT 1184.110 1676.780 1184.430 1676.840 ;
        RECT 1180.890 1676.640 1184.430 1676.780 ;
        RECT 1180.890 1676.580 1181.210 1676.640 ;
        RECT 1184.110 1676.580 1184.430 1676.640 ;
        RECT 341.390 19.620 341.710 19.680 ;
        RECT 1180.890 19.620 1181.210 19.680 ;
        RECT 341.390 19.480 1181.210 19.620 ;
        RECT 341.390 19.420 341.710 19.480 ;
        RECT 1180.890 19.420 1181.210 19.480 ;
      LAYER via ;
        RECT 1180.920 1676.580 1181.180 1676.840 ;
        RECT 1184.140 1676.580 1184.400 1676.840 ;
        RECT 341.420 19.420 341.680 19.680 ;
        RECT 1180.920 19.420 1181.180 19.680 ;
      LAYER met2 ;
        RECT 1184.500 1700.340 1184.780 1704.000 ;
        RECT 1184.500 1700.000 1184.800 1700.340 ;
        RECT 1184.660 1681.370 1184.800 1700.000 ;
        RECT 1184.200 1681.230 1184.800 1681.370 ;
        RECT 1184.200 1676.870 1184.340 1681.230 ;
        RECT 1180.920 1676.550 1181.180 1676.870 ;
        RECT 1184.140 1676.550 1184.400 1676.870 ;
        RECT 1180.980 19.710 1181.120 1676.550 ;
        RECT 341.420 19.390 341.680 19.710 ;
        RECT 1180.920 19.390 1181.180 19.710 ;
        RECT 341.480 2.400 341.620 19.390 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1181.350 1677.460 1181.670 1677.520 ;
        RECT 1186.410 1677.460 1186.730 1677.520 ;
        RECT 1181.350 1677.320 1186.730 1677.460 ;
        RECT 1181.350 1677.260 1181.670 1677.320 ;
        RECT 1186.410 1677.260 1186.730 1677.320 ;
        RECT 359.330 19.960 359.650 20.020 ;
        RECT 1181.350 19.960 1181.670 20.020 ;
        RECT 359.330 19.820 1181.670 19.960 ;
        RECT 359.330 19.760 359.650 19.820 ;
        RECT 1181.350 19.760 1181.670 19.820 ;
      LAYER via ;
        RECT 1181.380 1677.260 1181.640 1677.520 ;
        RECT 1186.440 1677.260 1186.700 1677.520 ;
        RECT 359.360 19.760 359.620 20.020 ;
        RECT 1181.380 19.760 1181.640 20.020 ;
      LAYER met2 ;
        RECT 1186.340 1700.340 1186.620 1704.000 ;
        RECT 1186.340 1700.000 1186.640 1700.340 ;
        RECT 1186.500 1677.550 1186.640 1700.000 ;
        RECT 1181.380 1677.230 1181.640 1677.550 ;
        RECT 1186.440 1677.230 1186.700 1677.550 ;
        RECT 1181.440 20.050 1181.580 1677.230 ;
        RECT 359.360 19.730 359.620 20.050 ;
        RECT 1181.380 19.730 1181.640 20.050 ;
        RECT 359.420 2.400 359.560 19.730 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1188.250 1678.480 1188.570 1678.540 ;
        RECT 1192.390 1678.480 1192.710 1678.540 ;
        RECT 1188.250 1678.340 1192.710 1678.480 ;
        RECT 1188.250 1678.280 1188.570 1678.340 ;
        RECT 1192.390 1678.280 1192.710 1678.340 ;
        RECT 420.510 20.300 420.830 20.360 ;
        RECT 1192.390 20.300 1192.710 20.360 ;
        RECT 420.510 20.160 1192.710 20.300 ;
        RECT 420.510 20.100 420.830 20.160 ;
        RECT 1192.390 20.100 1192.710 20.160 ;
        RECT 377.270 15.880 377.590 15.940 ;
        RECT 420.510 15.880 420.830 15.940 ;
        RECT 377.270 15.740 420.830 15.880 ;
        RECT 377.270 15.680 377.590 15.740 ;
        RECT 420.510 15.680 420.830 15.740 ;
      LAYER via ;
        RECT 1188.280 1678.280 1188.540 1678.540 ;
        RECT 1192.420 1678.280 1192.680 1678.540 ;
        RECT 420.540 20.100 420.800 20.360 ;
        RECT 1192.420 20.100 1192.680 20.360 ;
        RECT 377.300 15.680 377.560 15.940 ;
        RECT 420.540 15.680 420.800 15.940 ;
      LAYER met2 ;
        RECT 1188.180 1700.340 1188.460 1704.000 ;
        RECT 1188.180 1700.000 1188.480 1700.340 ;
        RECT 1188.340 1678.570 1188.480 1700.000 ;
        RECT 1188.280 1678.250 1188.540 1678.570 ;
        RECT 1192.420 1678.250 1192.680 1678.570 ;
        RECT 1192.480 20.390 1192.620 1678.250 ;
        RECT 420.540 20.070 420.800 20.390 ;
        RECT 1192.420 20.070 1192.680 20.390 ;
        RECT 420.600 15.970 420.740 20.070 ;
        RECT 377.300 15.650 377.560 15.970 ;
        RECT 420.540 15.650 420.800 15.970 ;
        RECT 377.360 2.400 377.500 15.650 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 395.210 20.640 395.530 20.700 ;
        RECT 1190.090 20.640 1190.410 20.700 ;
        RECT 395.210 20.500 1190.410 20.640 ;
        RECT 395.210 20.440 395.530 20.500 ;
        RECT 1190.090 20.440 1190.410 20.500 ;
      LAYER via ;
        RECT 395.240 20.440 395.500 20.700 ;
        RECT 1190.120 20.440 1190.380 20.700 ;
      LAYER met2 ;
        RECT 1190.020 1700.340 1190.300 1704.000 ;
        RECT 1190.020 1700.000 1190.320 1700.340 ;
        RECT 1190.180 20.730 1190.320 1700.000 ;
        RECT 395.240 20.410 395.500 20.730 ;
        RECT 1190.120 20.410 1190.380 20.730 ;
        RECT 395.300 2.400 395.440 20.410 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1125.305 16.235 1125.475 16.575 ;
        RECT 1125.305 16.065 1126.395 16.235 ;
      LAYER mcon ;
        RECT 1125.305 16.405 1125.475 16.575 ;
        RECT 1126.225 16.065 1126.395 16.235 ;
      LAYER met1 ;
        RECT 1190.550 1678.140 1190.870 1678.200 ;
        RECT 1191.930 1678.140 1192.250 1678.200 ;
        RECT 1190.550 1678.000 1192.250 1678.140 ;
        RECT 1190.550 1677.940 1190.870 1678.000 ;
        RECT 1191.930 1677.940 1192.250 1678.000 ;
        RECT 414.160 16.760 1125.460 16.900 ;
        RECT 413.150 16.220 413.470 16.280 ;
        RECT 414.160 16.220 414.300 16.760 ;
        RECT 1125.320 16.605 1125.460 16.760 ;
        RECT 1125.245 16.375 1125.535 16.605 ;
        RECT 413.150 16.080 414.300 16.220 ;
        RECT 1126.165 16.220 1126.455 16.265 ;
        RECT 1190.550 16.220 1190.870 16.280 ;
        RECT 1126.165 16.080 1190.870 16.220 ;
        RECT 413.150 16.020 413.470 16.080 ;
        RECT 1126.165 16.035 1126.455 16.080 ;
        RECT 1190.550 16.020 1190.870 16.080 ;
      LAYER via ;
        RECT 1190.580 1677.940 1190.840 1678.200 ;
        RECT 1191.960 1677.940 1192.220 1678.200 ;
        RECT 413.180 16.020 413.440 16.280 ;
        RECT 1190.580 16.020 1190.840 16.280 ;
      LAYER met2 ;
        RECT 1191.860 1700.340 1192.140 1704.000 ;
        RECT 1191.860 1700.000 1192.160 1700.340 ;
        RECT 1192.020 1678.230 1192.160 1700.000 ;
        RECT 1190.580 1677.910 1190.840 1678.230 ;
        RECT 1191.960 1677.910 1192.220 1678.230 ;
        RECT 1190.640 16.310 1190.780 1677.910 ;
        RECT 413.180 15.990 413.440 16.310 ;
        RECT 1190.580 15.990 1190.840 16.310 ;
        RECT 413.240 2.400 413.380 15.990 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.900 1700.340 1157.180 1704.000 ;
        RECT 1156.900 1700.000 1157.200 1700.340 ;
        RECT 1157.060 17.525 1157.200 1700.000 ;
        RECT 74.150 17.155 74.430 17.525 ;
        RECT 1156.990 17.155 1157.270 17.525 ;
        RECT 74.220 2.400 74.360 17.155 ;
        RECT 74.010 -4.800 74.570 2.400 ;
      LAYER via2 ;
        RECT 74.150 17.200 74.430 17.480 ;
        RECT 1156.990 17.200 1157.270 17.480 ;
      LAYER met3 ;
        RECT 74.125 17.490 74.455 17.505 ;
        RECT 1156.965 17.490 1157.295 17.505 ;
        RECT 74.125 17.190 1157.295 17.490 ;
        RECT 74.125 17.175 74.455 17.190 ;
        RECT 1156.965 17.175 1157.295 17.190 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1194.765 1159.145 1194.935 1207.255 ;
        RECT 1194.765 959.225 1194.935 1014.135 ;
        RECT 1124.845 16.745 1125.935 16.915 ;
        RECT 1124.845 16.405 1125.015 16.745 ;
        RECT 1145.545 13.685 1145.715 16.915 ;
        RECT 1170.845 13.685 1171.015 17.935 ;
      LAYER mcon ;
        RECT 1194.765 1207.085 1194.935 1207.255 ;
        RECT 1194.765 1013.965 1194.935 1014.135 ;
        RECT 1170.845 17.765 1171.015 17.935 ;
        RECT 1125.765 16.745 1125.935 16.915 ;
        RECT 1145.545 16.745 1145.715 16.915 ;
      LAYER met1 ;
        RECT 1194.230 1353.100 1194.550 1353.160 ;
        RECT 1194.230 1352.960 1194.920 1353.100 ;
        RECT 1194.230 1352.900 1194.550 1352.960 ;
        RECT 1194.780 1352.820 1194.920 1352.960 ;
        RECT 1194.690 1352.560 1195.010 1352.820 ;
        RECT 1194.690 1207.240 1195.010 1207.300 ;
        RECT 1194.495 1207.100 1195.010 1207.240 ;
        RECT 1194.690 1207.040 1195.010 1207.100 ;
        RECT 1194.690 1159.300 1195.010 1159.360 ;
        RECT 1194.495 1159.160 1195.010 1159.300 ;
        RECT 1194.690 1159.100 1195.010 1159.160 ;
        RECT 1194.690 1014.120 1195.010 1014.180 ;
        RECT 1194.495 1013.980 1195.010 1014.120 ;
        RECT 1194.690 1013.920 1195.010 1013.980 ;
        RECT 1194.690 959.380 1195.010 959.440 ;
        RECT 1194.495 959.240 1195.010 959.380 ;
        RECT 1194.690 959.180 1195.010 959.240 ;
        RECT 1193.770 814.200 1194.090 814.260 ;
        RECT 1194.690 814.200 1195.010 814.260 ;
        RECT 1193.770 814.060 1195.010 814.200 ;
        RECT 1193.770 814.000 1194.090 814.060 ;
        RECT 1194.690 814.000 1195.010 814.060 ;
        RECT 1170.785 17.920 1171.075 17.965 ;
        RECT 1194.690 17.920 1195.010 17.980 ;
        RECT 1170.785 17.780 1195.010 17.920 ;
        RECT 1170.785 17.735 1171.075 17.780 ;
        RECT 1194.690 17.720 1195.010 17.780 ;
        RECT 1125.705 16.900 1125.995 16.945 ;
        RECT 1145.485 16.900 1145.775 16.945 ;
        RECT 1125.705 16.760 1145.775 16.900 ;
        RECT 1125.705 16.715 1125.995 16.760 ;
        RECT 1145.485 16.715 1145.775 16.760 ;
        RECT 1124.785 16.560 1125.075 16.605 ;
        RECT 448.200 16.420 1125.075 16.560 ;
        RECT 430.630 16.220 430.950 16.280 ;
        RECT 448.200 16.220 448.340 16.420 ;
        RECT 1124.785 16.375 1125.075 16.420 ;
        RECT 430.630 16.080 448.340 16.220 ;
        RECT 430.630 16.020 430.950 16.080 ;
        RECT 1145.485 13.840 1145.775 13.885 ;
        RECT 1170.785 13.840 1171.075 13.885 ;
        RECT 1145.485 13.700 1171.075 13.840 ;
        RECT 1145.485 13.655 1145.775 13.700 ;
        RECT 1170.785 13.655 1171.075 13.700 ;
      LAYER via ;
        RECT 1194.260 1352.900 1194.520 1353.160 ;
        RECT 1194.720 1352.560 1194.980 1352.820 ;
        RECT 1194.720 1207.040 1194.980 1207.300 ;
        RECT 1194.720 1159.100 1194.980 1159.360 ;
        RECT 1194.720 1013.920 1194.980 1014.180 ;
        RECT 1194.720 959.180 1194.980 959.440 ;
        RECT 1193.800 814.000 1194.060 814.260 ;
        RECT 1194.720 814.000 1194.980 814.260 ;
        RECT 1194.720 17.720 1194.980 17.980 ;
        RECT 430.660 16.020 430.920 16.280 ;
      LAYER met2 ;
        RECT 1193.700 1700.410 1193.980 1704.000 ;
        RECT 1193.700 1700.270 1194.460 1700.410 ;
        RECT 1193.700 1700.000 1193.980 1700.270 ;
        RECT 1194.320 1669.130 1194.460 1700.270 ;
        RECT 1194.320 1668.990 1194.920 1669.130 ;
        RECT 1194.780 1400.530 1194.920 1668.990 ;
        RECT 1194.320 1400.390 1194.920 1400.530 ;
        RECT 1194.320 1353.190 1194.460 1400.390 ;
        RECT 1194.260 1352.870 1194.520 1353.190 ;
        RECT 1194.720 1352.530 1194.980 1352.850 ;
        RECT 1194.780 1207.330 1194.920 1352.530 ;
        RECT 1194.720 1207.010 1194.980 1207.330 ;
        RECT 1194.720 1159.070 1194.980 1159.390 ;
        RECT 1194.780 1014.210 1194.920 1159.070 ;
        RECT 1194.720 1013.890 1194.980 1014.210 ;
        RECT 1194.720 959.150 1194.980 959.470 ;
        RECT 1194.780 814.290 1194.920 959.150 ;
        RECT 1193.800 813.970 1194.060 814.290 ;
        RECT 1194.720 813.970 1194.980 814.290 ;
        RECT 1193.860 766.205 1194.000 813.970 ;
        RECT 1193.790 765.835 1194.070 766.205 ;
        RECT 1194.710 765.835 1194.990 766.205 ;
        RECT 1194.780 725.405 1194.920 765.835 ;
        RECT 1194.710 725.035 1194.990 725.405 ;
        RECT 1193.790 723.675 1194.070 724.045 ;
        RECT 1193.860 676.445 1194.000 723.675 ;
        RECT 1193.790 676.075 1194.070 676.445 ;
        RECT 1194.710 676.075 1194.990 676.445 ;
        RECT 1194.780 628.845 1194.920 676.075 ;
        RECT 1194.710 628.475 1194.990 628.845 ;
        RECT 1193.790 626.435 1194.070 626.805 ;
        RECT 1193.860 579.885 1194.000 626.435 ;
        RECT 1193.790 579.515 1194.070 579.885 ;
        RECT 1194.710 579.515 1194.990 579.885 ;
        RECT 1194.780 18.010 1194.920 579.515 ;
        RECT 1194.720 17.690 1194.980 18.010 ;
        RECT 430.660 15.990 430.920 16.310 ;
        RECT 430.720 2.400 430.860 15.990 ;
        RECT 430.510 -4.800 431.070 2.400 ;
      LAYER via2 ;
        RECT 1193.790 765.880 1194.070 766.160 ;
        RECT 1194.710 765.880 1194.990 766.160 ;
        RECT 1194.710 725.080 1194.990 725.360 ;
        RECT 1193.790 723.720 1194.070 724.000 ;
        RECT 1193.790 676.120 1194.070 676.400 ;
        RECT 1194.710 676.120 1194.990 676.400 ;
        RECT 1194.710 628.520 1194.990 628.800 ;
        RECT 1193.790 626.480 1194.070 626.760 ;
        RECT 1193.790 579.560 1194.070 579.840 ;
        RECT 1194.710 579.560 1194.990 579.840 ;
      LAYER met3 ;
        RECT 1193.765 766.170 1194.095 766.185 ;
        RECT 1194.685 766.170 1195.015 766.185 ;
        RECT 1193.765 765.870 1195.015 766.170 ;
        RECT 1193.765 765.855 1194.095 765.870 ;
        RECT 1194.685 765.855 1195.015 765.870 ;
        RECT 1194.685 725.370 1195.015 725.385 ;
        RECT 1194.470 725.055 1195.015 725.370 ;
        RECT 1193.765 724.010 1194.095 724.025 ;
        RECT 1194.470 724.010 1194.770 725.055 ;
        RECT 1193.765 723.710 1194.770 724.010 ;
        RECT 1193.765 723.695 1194.095 723.710 ;
        RECT 1193.765 676.410 1194.095 676.425 ;
        RECT 1194.685 676.410 1195.015 676.425 ;
        RECT 1193.765 676.110 1195.015 676.410 ;
        RECT 1193.765 676.095 1194.095 676.110 ;
        RECT 1194.685 676.095 1195.015 676.110 ;
        RECT 1194.685 628.810 1195.015 628.825 ;
        RECT 1194.470 628.495 1195.015 628.810 ;
        RECT 1193.765 626.770 1194.095 626.785 ;
        RECT 1194.470 626.770 1194.770 628.495 ;
        RECT 1193.765 626.470 1194.770 626.770 ;
        RECT 1193.765 626.455 1194.095 626.470 ;
        RECT 1193.765 579.850 1194.095 579.865 ;
        RECT 1194.685 579.850 1195.015 579.865 ;
        RECT 1193.765 579.550 1195.015 579.850 ;
        RECT 1193.765 579.535 1194.095 579.550 ;
        RECT 1194.685 579.535 1195.015 579.550 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1148.765 15.045 1148.935 16.575 ;
      LAYER mcon ;
        RECT 1148.765 16.405 1148.935 16.575 ;
      LAYER met1 ;
        RECT 1195.610 1678.480 1195.930 1678.540 ;
        RECT 1199.750 1678.480 1200.070 1678.540 ;
        RECT 1195.610 1678.340 1200.070 1678.480 ;
        RECT 1195.610 1678.280 1195.930 1678.340 ;
        RECT 1199.750 1678.280 1200.070 1678.340 ;
        RECT 1148.705 16.560 1148.995 16.605 ;
        RECT 1125.780 16.420 1148.995 16.560 ;
        RECT 448.570 16.220 448.890 16.280 ;
        RECT 1125.780 16.220 1125.920 16.420 ;
        RECT 1148.705 16.375 1148.995 16.420 ;
        RECT 448.570 16.080 1125.920 16.220 ;
        RECT 448.570 16.020 448.890 16.080 ;
        RECT 1148.705 15.200 1148.995 15.245 ;
        RECT 1199.750 15.200 1200.070 15.260 ;
        RECT 1148.705 15.060 1200.070 15.200 ;
        RECT 1148.705 15.015 1148.995 15.060 ;
        RECT 1199.750 15.000 1200.070 15.060 ;
      LAYER via ;
        RECT 1195.640 1678.280 1195.900 1678.540 ;
        RECT 1199.780 1678.280 1200.040 1678.540 ;
        RECT 448.600 16.020 448.860 16.280 ;
        RECT 1199.780 15.000 1200.040 15.260 ;
      LAYER met2 ;
        RECT 1195.540 1700.340 1195.820 1704.000 ;
        RECT 1195.540 1700.000 1195.840 1700.340 ;
        RECT 1195.700 1678.570 1195.840 1700.000 ;
        RECT 1195.640 1678.250 1195.900 1678.570 ;
        RECT 1199.780 1678.250 1200.040 1678.570 ;
        RECT 448.600 15.990 448.860 16.310 ;
        RECT 448.660 2.400 448.800 15.990 ;
        RECT 1199.840 15.290 1199.980 1678.250 ;
        RECT 1199.780 14.970 1200.040 15.290 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 466.510 15.880 466.830 15.940 ;
        RECT 1197.450 15.880 1197.770 15.940 ;
        RECT 466.510 15.740 1197.770 15.880 ;
        RECT 466.510 15.680 466.830 15.740 ;
        RECT 1197.450 15.680 1197.770 15.740 ;
      LAYER via ;
        RECT 466.540 15.680 466.800 15.940 ;
        RECT 1197.480 15.680 1197.740 15.940 ;
      LAYER met2 ;
        RECT 1197.380 1700.340 1197.660 1704.000 ;
        RECT 1197.380 1700.000 1197.680 1700.340 ;
        RECT 1197.540 15.970 1197.680 1700.000 ;
        RECT 466.540 15.650 466.800 15.970 ;
        RECT 1197.480 15.650 1197.740 15.970 ;
        RECT 466.600 2.400 466.740 15.650 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1197.910 1678.140 1198.230 1678.200 ;
        RECT 1199.290 1678.140 1199.610 1678.200 ;
        RECT 1197.910 1678.000 1199.610 1678.140 ;
        RECT 1197.910 1677.940 1198.230 1678.000 ;
        RECT 1199.290 1677.940 1199.610 1678.000 ;
        RECT 1198.370 15.540 1198.690 15.600 ;
        RECT 541.580 15.400 1198.690 15.540 ;
        RECT 484.450 15.200 484.770 15.260 ;
        RECT 541.580 15.200 541.720 15.400 ;
        RECT 1198.370 15.340 1198.690 15.400 ;
        RECT 484.450 15.060 541.720 15.200 ;
        RECT 484.450 15.000 484.770 15.060 ;
      LAYER via ;
        RECT 1197.940 1677.940 1198.200 1678.200 ;
        RECT 1199.320 1677.940 1199.580 1678.200 ;
        RECT 484.480 15.000 484.740 15.260 ;
        RECT 1198.400 15.340 1198.660 15.600 ;
      LAYER met2 ;
        RECT 1199.220 1700.340 1199.500 1704.000 ;
        RECT 1199.220 1700.000 1199.520 1700.340 ;
        RECT 1199.380 1678.230 1199.520 1700.000 ;
        RECT 1197.940 1677.910 1198.200 1678.230 ;
        RECT 1199.320 1677.910 1199.580 1678.230 ;
        RECT 1198.000 21.490 1198.140 1677.910 ;
        RECT 1198.000 21.350 1198.600 21.490 ;
        RECT 1198.460 15.630 1198.600 21.350 ;
        RECT 1198.400 15.310 1198.660 15.630 ;
        RECT 484.480 14.970 484.740 15.290 ;
        RECT 484.540 2.400 484.680 14.970 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1201.130 1689.840 1201.450 1690.100 ;
        RECT 1201.220 1689.700 1201.360 1689.840 ;
        RECT 1186.960 1689.560 1201.360 1689.700 ;
        RECT 503.310 1689.360 503.630 1689.420 ;
        RECT 1186.960 1689.360 1187.100 1689.560 ;
        RECT 503.310 1689.220 1187.100 1689.360 ;
        RECT 503.310 1689.160 503.630 1689.220 ;
      LAYER via ;
        RECT 1201.160 1689.840 1201.420 1690.100 ;
        RECT 503.340 1689.160 503.600 1689.420 ;
      LAYER met2 ;
        RECT 1201.060 1700.340 1201.340 1704.000 ;
        RECT 1201.060 1700.000 1201.360 1700.340 ;
        RECT 1201.220 1690.130 1201.360 1700.000 ;
        RECT 1201.160 1689.810 1201.420 1690.130 ;
        RECT 503.340 1689.130 503.600 1689.450 ;
        RECT 503.400 24.210 503.540 1689.130 ;
        RECT 502.480 24.070 503.540 24.210 ;
        RECT 502.480 2.400 502.620 24.070 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1203.430 1678.140 1203.750 1678.200 ;
        RECT 1205.270 1678.140 1205.590 1678.200 ;
        RECT 1203.430 1678.000 1205.590 1678.140 ;
        RECT 1203.430 1677.940 1203.750 1678.000 ;
        RECT 1205.270 1677.940 1205.590 1678.000 ;
        RECT 542.040 15.060 1131.900 15.200 ;
        RECT 519.870 14.520 520.190 14.580 ;
        RECT 542.040 14.520 542.180 15.060 ;
        RECT 1131.760 14.860 1131.900 15.060 ;
        RECT 1205.270 14.860 1205.590 14.920 ;
        RECT 1131.760 14.720 1205.590 14.860 ;
        RECT 1205.270 14.660 1205.590 14.720 ;
        RECT 519.870 14.380 542.180 14.520 ;
        RECT 519.870 14.320 520.190 14.380 ;
      LAYER via ;
        RECT 1203.460 1677.940 1203.720 1678.200 ;
        RECT 1205.300 1677.940 1205.560 1678.200 ;
        RECT 519.900 14.320 520.160 14.580 ;
        RECT 1205.300 14.660 1205.560 14.920 ;
      LAYER met2 ;
        RECT 1202.900 1700.410 1203.180 1704.000 ;
        RECT 1202.900 1700.270 1203.660 1700.410 ;
        RECT 1202.900 1700.000 1203.180 1700.270 ;
        RECT 1203.520 1678.230 1203.660 1700.270 ;
        RECT 1203.460 1677.910 1203.720 1678.230 ;
        RECT 1205.300 1677.910 1205.560 1678.230 ;
        RECT 1205.360 14.950 1205.500 1677.910 ;
        RECT 1205.300 14.630 1205.560 14.950 ;
        RECT 519.900 14.290 520.160 14.610 ;
        RECT 519.960 2.400 520.100 14.290 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1204.810 1690.380 1205.130 1690.440 ;
        RECT 1188.800 1690.240 1205.130 1690.380 ;
        RECT 537.810 1690.040 538.130 1690.100 ;
        RECT 1188.800 1690.040 1188.940 1690.240 ;
        RECT 1204.810 1690.180 1205.130 1690.240 ;
        RECT 537.810 1689.900 1188.940 1690.040 ;
        RECT 537.810 1689.840 538.130 1689.900 ;
      LAYER via ;
        RECT 537.840 1689.840 538.100 1690.100 ;
        RECT 1204.840 1690.180 1205.100 1690.440 ;
      LAYER met2 ;
        RECT 1204.740 1700.340 1205.020 1704.000 ;
        RECT 1204.740 1700.000 1205.040 1700.340 ;
        RECT 1204.900 1690.470 1205.040 1700.000 ;
        RECT 1204.840 1690.150 1205.100 1690.470 ;
        RECT 537.840 1689.810 538.100 1690.130 ;
        RECT 537.900 2.400 538.040 1689.810 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1131.285 14.705 1131.455 17.935 ;
        RECT 1149.225 17.765 1149.395 18.615 ;
      LAYER mcon ;
        RECT 1149.225 18.445 1149.395 18.615 ;
        RECT 1131.285 17.765 1131.455 17.935 ;
      LAYER met1 ;
        RECT 1149.165 18.600 1149.455 18.645 ;
        RECT 1206.650 18.600 1206.970 18.660 ;
        RECT 1149.165 18.460 1206.970 18.600 ;
        RECT 1149.165 18.415 1149.455 18.460 ;
        RECT 1206.650 18.400 1206.970 18.460 ;
        RECT 1131.225 17.920 1131.515 17.965 ;
        RECT 1149.165 17.920 1149.455 17.965 ;
        RECT 1131.225 17.780 1149.455 17.920 ;
        RECT 1131.225 17.735 1131.515 17.780 ;
        RECT 1149.165 17.735 1149.455 17.780 ;
        RECT 1131.225 14.860 1131.515 14.905 ;
        RECT 572.860 14.720 1131.515 14.860 ;
        RECT 555.750 14.520 556.070 14.580 ;
        RECT 572.860 14.520 573.000 14.720 ;
        RECT 1131.225 14.675 1131.515 14.720 ;
        RECT 555.750 14.380 573.000 14.520 ;
        RECT 555.750 14.320 556.070 14.380 ;
      LAYER via ;
        RECT 1206.680 18.400 1206.940 18.660 ;
        RECT 555.780 14.320 556.040 14.580 ;
      LAYER met2 ;
        RECT 1206.580 1700.340 1206.860 1704.000 ;
        RECT 1206.580 1700.000 1206.880 1700.340 ;
        RECT 1206.740 18.690 1206.880 1700.000 ;
        RECT 1206.680 18.370 1206.940 18.690 ;
        RECT 555.780 14.290 556.040 14.610 ;
        RECT 555.840 2.400 555.980 14.290 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1186.485 1688.865 1186.655 1689.715 ;
      LAYER mcon ;
        RECT 1186.485 1689.545 1186.655 1689.715 ;
      LAYER met1 ;
        RECT 579.210 1689.700 579.530 1689.760 ;
        RECT 1186.425 1689.700 1186.715 1689.745 ;
        RECT 579.210 1689.560 1186.715 1689.700 ;
        RECT 579.210 1689.500 579.530 1689.560 ;
        RECT 1186.425 1689.515 1186.715 1689.560 ;
        RECT 1186.425 1689.020 1186.715 1689.065 ;
        RECT 1208.490 1689.020 1208.810 1689.080 ;
        RECT 1186.425 1688.880 1208.810 1689.020 ;
        RECT 1186.425 1688.835 1186.715 1688.880 ;
        RECT 1208.490 1688.820 1208.810 1688.880 ;
        RECT 573.690 14.520 574.010 14.580 ;
        RECT 579.210 14.520 579.530 14.580 ;
        RECT 573.690 14.380 579.530 14.520 ;
        RECT 573.690 14.320 574.010 14.380 ;
        RECT 579.210 14.320 579.530 14.380 ;
      LAYER via ;
        RECT 579.240 1689.500 579.500 1689.760 ;
        RECT 1208.520 1688.820 1208.780 1689.080 ;
        RECT 573.720 14.320 573.980 14.580 ;
        RECT 579.240 14.320 579.500 14.580 ;
      LAYER met2 ;
        RECT 1208.420 1700.340 1208.700 1704.000 ;
        RECT 1208.420 1700.000 1208.720 1700.340 ;
        RECT 579.240 1689.470 579.500 1689.790 ;
        RECT 579.300 14.610 579.440 1689.470 ;
        RECT 1208.580 1689.110 1208.720 1700.000 ;
        RECT 1208.520 1688.790 1208.780 1689.110 ;
        RECT 573.720 14.290 573.980 14.610 ;
        RECT 579.240 14.290 579.500 14.610 ;
        RECT 573.780 2.400 573.920 14.290 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1210.330 14.520 1210.650 14.580 ;
        RECT 607.360 14.380 1210.650 14.520 ;
        RECT 591.170 14.180 591.490 14.240 ;
        RECT 607.360 14.180 607.500 14.380 ;
        RECT 1210.330 14.320 1210.650 14.380 ;
        RECT 591.170 14.040 607.500 14.180 ;
        RECT 591.170 13.980 591.490 14.040 ;
      LAYER via ;
        RECT 591.200 13.980 591.460 14.240 ;
        RECT 1210.360 14.320 1210.620 14.580 ;
      LAYER met2 ;
        RECT 1210.260 1700.340 1210.540 1704.000 ;
        RECT 1210.260 1700.000 1210.560 1700.340 ;
        RECT 1210.420 14.610 1210.560 1700.000 ;
        RECT 1210.360 14.290 1210.620 14.610 ;
        RECT 591.200 13.950 591.460 14.270 ;
        RECT 591.260 2.400 591.400 13.950 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 161.990 1688.340 162.310 1688.400 ;
        RECT 1159.730 1688.340 1160.050 1688.400 ;
        RECT 161.990 1688.200 1160.050 1688.340 ;
        RECT 161.990 1688.140 162.310 1688.200 ;
        RECT 1159.730 1688.140 1160.050 1688.200 ;
        RECT 161.990 17.580 162.310 17.640 ;
        RECT 143.680 17.440 162.310 17.580 ;
        RECT 97.590 17.240 97.910 17.300 ;
        RECT 143.680 17.240 143.820 17.440 ;
        RECT 161.990 17.380 162.310 17.440 ;
        RECT 97.590 17.100 143.820 17.240 ;
        RECT 97.590 17.040 97.910 17.100 ;
      LAYER via ;
        RECT 162.020 1688.140 162.280 1688.400 ;
        RECT 1159.760 1688.140 1160.020 1688.400 ;
        RECT 97.620 17.040 97.880 17.300 ;
        RECT 162.020 17.380 162.280 17.640 ;
      LAYER met2 ;
        RECT 1159.660 1700.340 1159.940 1704.000 ;
        RECT 1159.660 1700.000 1159.960 1700.340 ;
        RECT 1159.820 1688.430 1159.960 1700.000 ;
        RECT 162.020 1688.110 162.280 1688.430 ;
        RECT 1159.760 1688.110 1160.020 1688.430 ;
        RECT 162.080 17.670 162.220 1688.110 ;
        RECT 162.020 17.350 162.280 17.670 ;
        RECT 97.620 17.010 97.880 17.330 ;
        RECT 97.680 2.400 97.820 17.010 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1210.790 1678.140 1211.110 1678.200 ;
        RECT 1212.170 1678.140 1212.490 1678.200 ;
        RECT 1210.790 1678.000 1212.490 1678.140 ;
        RECT 1210.790 1677.940 1211.110 1678.000 ;
        RECT 1212.170 1677.940 1212.490 1678.000 ;
        RECT 609.110 14.180 609.430 14.240 ;
        RECT 1210.790 14.180 1211.110 14.240 ;
        RECT 609.110 14.040 1211.110 14.180 ;
        RECT 609.110 13.980 609.430 14.040 ;
        RECT 1210.790 13.980 1211.110 14.040 ;
      LAYER via ;
        RECT 1210.820 1677.940 1211.080 1678.200 ;
        RECT 1212.200 1677.940 1212.460 1678.200 ;
        RECT 609.140 13.980 609.400 14.240 ;
        RECT 1210.820 13.980 1211.080 14.240 ;
      LAYER met2 ;
        RECT 1212.100 1700.340 1212.380 1704.000 ;
        RECT 1212.100 1700.000 1212.400 1700.340 ;
        RECT 1212.260 1678.230 1212.400 1700.000 ;
        RECT 1210.820 1677.910 1211.080 1678.230 ;
        RECT 1212.200 1677.910 1212.460 1678.230 ;
        RECT 1210.880 14.270 1211.020 1677.910 ;
        RECT 609.140 13.950 609.400 14.270 ;
        RECT 1210.820 13.950 1211.080 14.270 ;
        RECT 609.200 2.400 609.340 13.950 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1188.325 1688.525 1188.495 1690.395 ;
      LAYER mcon ;
        RECT 1188.325 1690.225 1188.495 1690.395 ;
      LAYER met1 ;
        RECT 627.510 1690.380 627.830 1690.440 ;
        RECT 1188.265 1690.380 1188.555 1690.425 ;
        RECT 627.510 1690.240 1188.555 1690.380 ;
        RECT 627.510 1690.180 627.830 1690.240 ;
        RECT 1188.265 1690.195 1188.555 1690.240 ;
        RECT 1188.265 1688.680 1188.555 1688.725 ;
        RECT 1214.010 1688.680 1214.330 1688.740 ;
        RECT 1188.265 1688.540 1214.330 1688.680 ;
        RECT 1188.265 1688.495 1188.555 1688.540 ;
        RECT 1214.010 1688.480 1214.330 1688.540 ;
      LAYER via ;
        RECT 627.540 1690.180 627.800 1690.440 ;
        RECT 1214.040 1688.480 1214.300 1688.740 ;
      LAYER met2 ;
        RECT 1213.940 1700.340 1214.220 1704.000 ;
        RECT 1213.940 1700.000 1214.240 1700.340 ;
        RECT 627.540 1690.150 627.800 1690.470 ;
        RECT 627.600 17.410 627.740 1690.150 ;
        RECT 1214.100 1688.770 1214.240 1700.000 ;
        RECT 1214.040 1688.450 1214.300 1688.770 ;
        RECT 627.140 17.270 627.740 17.410 ;
        RECT 627.140 2.400 627.280 17.270 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1161.570 1678.140 1161.890 1678.200 ;
        RECT 1163.870 1678.140 1164.190 1678.200 ;
        RECT 1161.570 1678.000 1164.190 1678.140 ;
        RECT 1161.570 1677.940 1161.890 1678.000 ;
        RECT 1163.870 1677.940 1164.190 1678.000 ;
      LAYER via ;
        RECT 1161.600 1677.940 1161.860 1678.200 ;
        RECT 1163.900 1677.940 1164.160 1678.200 ;
      LAYER met2 ;
        RECT 1161.960 1700.340 1162.240 1704.000 ;
        RECT 1161.960 1700.000 1162.260 1700.340 ;
        RECT 1162.120 1699.730 1162.260 1700.000 ;
        RECT 1161.660 1699.590 1162.260 1699.730 ;
        RECT 1161.660 1678.230 1161.800 1699.590 ;
        RECT 1161.600 1677.910 1161.860 1678.230 ;
        RECT 1163.900 1677.910 1164.160 1678.230 ;
        RECT 1163.960 18.885 1164.100 1677.910 ;
        RECT 121.530 18.515 121.810 18.885 ;
        RECT 1163.890 18.515 1164.170 18.885 ;
        RECT 121.600 2.400 121.740 18.515 ;
        RECT 121.390 -4.800 121.950 2.400 ;
      LAYER via2 ;
        RECT 121.530 18.560 121.810 18.840 ;
        RECT 1163.890 18.560 1164.170 18.840 ;
      LAYER met3 ;
        RECT 121.505 18.850 121.835 18.865 ;
        RECT 1163.865 18.850 1164.195 18.865 ;
        RECT 121.505 18.550 1164.195 18.850 ;
        RECT 121.505 18.535 121.835 18.550 ;
        RECT 1163.865 18.535 1164.195 18.550 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 175.790 1689.020 176.110 1689.080 ;
        RECT 1164.330 1689.020 1164.650 1689.080 ;
        RECT 175.790 1688.880 1164.650 1689.020 ;
        RECT 175.790 1688.820 176.110 1688.880 ;
        RECT 1164.330 1688.820 1164.650 1688.880 ;
        RECT 145.430 17.240 145.750 17.300 ;
        RECT 175.790 17.240 176.110 17.300 ;
        RECT 145.430 17.100 176.110 17.240 ;
        RECT 145.430 17.040 145.750 17.100 ;
        RECT 175.790 17.040 176.110 17.100 ;
      LAYER via ;
        RECT 175.820 1688.820 176.080 1689.080 ;
        RECT 1164.360 1688.820 1164.620 1689.080 ;
        RECT 145.460 17.040 145.720 17.300 ;
        RECT 175.820 17.040 176.080 17.300 ;
      LAYER met2 ;
        RECT 1164.260 1700.340 1164.540 1704.000 ;
        RECT 1164.260 1700.000 1164.560 1700.340 ;
        RECT 1164.420 1689.110 1164.560 1700.000 ;
        RECT 175.820 1688.790 176.080 1689.110 ;
        RECT 1164.360 1688.790 1164.620 1689.110 ;
        RECT 175.880 17.330 176.020 1688.790 ;
        RECT 145.460 17.010 145.720 17.330 ;
        RECT 175.820 17.010 176.080 17.330 ;
        RECT 145.520 2.400 145.660 17.010 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1169.925 1635.485 1170.095 1671.695 ;
        RECT 1169.005 476.085 1169.175 524.195 ;
      LAYER mcon ;
        RECT 1169.925 1671.525 1170.095 1671.695 ;
        RECT 1169.005 524.025 1169.175 524.195 ;
      LAYER met1 ;
        RECT 1166.630 1671.680 1166.950 1671.740 ;
        RECT 1169.865 1671.680 1170.155 1671.725 ;
        RECT 1166.630 1671.540 1170.155 1671.680 ;
        RECT 1166.630 1671.480 1166.950 1671.540 ;
        RECT 1169.865 1671.495 1170.155 1671.540 ;
        RECT 1169.850 1635.640 1170.170 1635.700 ;
        RECT 1169.655 1635.500 1170.170 1635.640 ;
        RECT 1169.850 1635.440 1170.170 1635.500 ;
        RECT 1169.850 1594.300 1170.170 1594.560 ;
        RECT 1169.940 1593.880 1170.080 1594.300 ;
        RECT 1169.850 1593.620 1170.170 1593.880 ;
        RECT 1169.850 1538.540 1170.170 1538.800 ;
        RECT 1168.930 1538.400 1169.250 1538.460 ;
        RECT 1169.940 1538.400 1170.080 1538.540 ;
        RECT 1168.930 1538.260 1170.080 1538.400 ;
        RECT 1168.930 1538.200 1169.250 1538.260 ;
        RECT 1168.470 1414.640 1168.790 1414.700 ;
        RECT 1169.390 1414.640 1169.710 1414.700 ;
        RECT 1168.470 1414.500 1169.710 1414.640 ;
        RECT 1168.470 1414.440 1168.790 1414.500 ;
        RECT 1169.390 1414.440 1169.710 1414.500 ;
        RECT 1168.470 1318.080 1168.790 1318.140 ;
        RECT 1169.390 1318.080 1169.710 1318.140 ;
        RECT 1168.470 1317.940 1169.710 1318.080 ;
        RECT 1168.470 1317.880 1168.790 1317.940 ;
        RECT 1169.390 1317.880 1169.710 1317.940 ;
        RECT 1168.470 1221.520 1168.790 1221.580 ;
        RECT 1169.390 1221.520 1169.710 1221.580 ;
        RECT 1168.470 1221.380 1169.710 1221.520 ;
        RECT 1168.470 1221.320 1168.790 1221.380 ;
        RECT 1169.390 1221.320 1169.710 1221.380 ;
        RECT 1168.470 1124.960 1168.790 1125.020 ;
        RECT 1169.390 1124.960 1169.710 1125.020 ;
        RECT 1168.470 1124.820 1169.710 1124.960 ;
        RECT 1168.470 1124.760 1168.790 1124.820 ;
        RECT 1169.390 1124.760 1169.710 1124.820 ;
        RECT 1168.470 1028.400 1168.790 1028.460 ;
        RECT 1169.390 1028.400 1169.710 1028.460 ;
        RECT 1168.470 1028.260 1169.710 1028.400 ;
        RECT 1168.470 1028.200 1168.790 1028.260 ;
        RECT 1169.390 1028.200 1169.710 1028.260 ;
        RECT 1168.470 931.840 1168.790 931.900 ;
        RECT 1169.390 931.840 1169.710 931.900 ;
        RECT 1168.470 931.700 1169.710 931.840 ;
        RECT 1168.470 931.640 1168.790 931.700 ;
        RECT 1169.390 931.640 1169.710 931.700 ;
        RECT 1168.470 835.280 1168.790 835.340 ;
        RECT 1169.390 835.280 1169.710 835.340 ;
        RECT 1168.470 835.140 1169.710 835.280 ;
        RECT 1168.470 835.080 1168.790 835.140 ;
        RECT 1169.390 835.080 1169.710 835.140 ;
        RECT 1168.470 641.820 1168.790 641.880 ;
        RECT 1169.390 641.820 1169.710 641.880 ;
        RECT 1168.470 641.680 1169.710 641.820 ;
        RECT 1168.470 641.620 1168.790 641.680 ;
        RECT 1169.390 641.620 1169.710 641.680 ;
        RECT 1168.470 545.260 1168.790 545.320 ;
        RECT 1169.390 545.260 1169.710 545.320 ;
        RECT 1168.470 545.120 1169.710 545.260 ;
        RECT 1168.470 545.060 1168.790 545.120 ;
        RECT 1169.390 545.060 1169.710 545.120 ;
        RECT 1168.930 524.180 1169.250 524.240 ;
        RECT 1168.735 524.040 1169.250 524.180 ;
        RECT 1168.930 523.980 1169.250 524.040 ;
        RECT 1168.945 476.240 1169.235 476.285 ;
        RECT 1169.850 476.240 1170.170 476.300 ;
        RECT 1168.945 476.100 1170.170 476.240 ;
        RECT 1168.945 476.055 1169.235 476.100 ;
        RECT 1169.850 476.040 1170.170 476.100 ;
        RECT 1168.930 386.480 1169.250 386.540 ;
        RECT 1169.390 386.480 1169.710 386.540 ;
        RECT 1168.930 386.340 1169.710 386.480 ;
        RECT 1168.930 386.280 1169.250 386.340 ;
        RECT 1169.390 386.280 1169.710 386.340 ;
        RECT 1168.930 338.200 1169.250 338.260 ;
        RECT 1169.390 338.200 1169.710 338.260 ;
        RECT 1168.930 338.060 1169.710 338.200 ;
        RECT 1168.930 338.000 1169.250 338.060 ;
        RECT 1169.390 338.000 1169.710 338.060 ;
      LAYER via ;
        RECT 1166.660 1671.480 1166.920 1671.740 ;
        RECT 1169.880 1635.440 1170.140 1635.700 ;
        RECT 1169.880 1594.300 1170.140 1594.560 ;
        RECT 1169.880 1593.620 1170.140 1593.880 ;
        RECT 1169.880 1538.540 1170.140 1538.800 ;
        RECT 1168.960 1538.200 1169.220 1538.460 ;
        RECT 1168.500 1414.440 1168.760 1414.700 ;
        RECT 1169.420 1414.440 1169.680 1414.700 ;
        RECT 1168.500 1317.880 1168.760 1318.140 ;
        RECT 1169.420 1317.880 1169.680 1318.140 ;
        RECT 1168.500 1221.320 1168.760 1221.580 ;
        RECT 1169.420 1221.320 1169.680 1221.580 ;
        RECT 1168.500 1124.760 1168.760 1125.020 ;
        RECT 1169.420 1124.760 1169.680 1125.020 ;
        RECT 1168.500 1028.200 1168.760 1028.460 ;
        RECT 1169.420 1028.200 1169.680 1028.460 ;
        RECT 1168.500 931.640 1168.760 931.900 ;
        RECT 1169.420 931.640 1169.680 931.900 ;
        RECT 1168.500 835.080 1168.760 835.340 ;
        RECT 1169.420 835.080 1169.680 835.340 ;
        RECT 1168.500 641.620 1168.760 641.880 ;
        RECT 1169.420 641.620 1169.680 641.880 ;
        RECT 1168.500 545.060 1168.760 545.320 ;
        RECT 1169.420 545.060 1169.680 545.320 ;
        RECT 1168.960 523.980 1169.220 524.240 ;
        RECT 1169.880 476.040 1170.140 476.300 ;
        RECT 1168.960 386.280 1169.220 386.540 ;
        RECT 1169.420 386.280 1169.680 386.540 ;
        RECT 1168.960 338.000 1169.220 338.260 ;
        RECT 1169.420 338.000 1169.680 338.260 ;
      LAYER met2 ;
        RECT 1166.100 1700.410 1166.380 1704.000 ;
        RECT 1166.100 1700.270 1166.860 1700.410 ;
        RECT 1166.100 1700.000 1166.380 1700.270 ;
        RECT 1166.720 1671.770 1166.860 1700.270 ;
        RECT 1166.660 1671.450 1166.920 1671.770 ;
        RECT 1169.880 1635.410 1170.140 1635.730 ;
        RECT 1169.940 1594.590 1170.080 1635.410 ;
        RECT 1169.880 1594.270 1170.140 1594.590 ;
        RECT 1169.880 1593.590 1170.140 1593.910 ;
        RECT 1169.940 1538.830 1170.080 1593.590 ;
        RECT 1169.880 1538.510 1170.140 1538.830 ;
        RECT 1168.960 1538.170 1169.220 1538.490 ;
        RECT 1169.020 1473.290 1169.160 1538.170 ;
        RECT 1169.020 1473.150 1169.620 1473.290 ;
        RECT 1169.480 1414.730 1169.620 1473.150 ;
        RECT 1168.500 1414.410 1168.760 1414.730 ;
        RECT 1169.420 1414.410 1169.680 1414.730 ;
        RECT 1168.560 1414.130 1168.700 1414.410 ;
        RECT 1168.560 1413.990 1169.160 1414.130 ;
        RECT 1169.020 1366.530 1169.160 1413.990 ;
        RECT 1169.020 1366.390 1169.620 1366.530 ;
        RECT 1169.480 1318.170 1169.620 1366.390 ;
        RECT 1168.500 1317.850 1168.760 1318.170 ;
        RECT 1169.420 1317.850 1169.680 1318.170 ;
        RECT 1168.560 1317.570 1168.700 1317.850 ;
        RECT 1168.560 1317.430 1169.160 1317.570 ;
        RECT 1169.020 1269.970 1169.160 1317.430 ;
        RECT 1169.020 1269.830 1169.620 1269.970 ;
        RECT 1169.480 1221.610 1169.620 1269.830 ;
        RECT 1168.500 1221.290 1168.760 1221.610 ;
        RECT 1169.420 1221.290 1169.680 1221.610 ;
        RECT 1168.560 1221.010 1168.700 1221.290 ;
        RECT 1168.560 1220.870 1169.160 1221.010 ;
        RECT 1169.020 1173.410 1169.160 1220.870 ;
        RECT 1169.020 1173.270 1169.620 1173.410 ;
        RECT 1169.480 1125.050 1169.620 1173.270 ;
        RECT 1168.500 1124.730 1168.760 1125.050 ;
        RECT 1169.420 1124.730 1169.680 1125.050 ;
        RECT 1168.560 1124.450 1168.700 1124.730 ;
        RECT 1168.560 1124.310 1169.160 1124.450 ;
        RECT 1169.020 1076.850 1169.160 1124.310 ;
        RECT 1169.020 1076.710 1169.620 1076.850 ;
        RECT 1169.480 1028.490 1169.620 1076.710 ;
        RECT 1168.500 1028.170 1168.760 1028.490 ;
        RECT 1169.420 1028.170 1169.680 1028.490 ;
        RECT 1168.560 1027.890 1168.700 1028.170 ;
        RECT 1168.560 1027.750 1169.160 1027.890 ;
        RECT 1169.020 980.290 1169.160 1027.750 ;
        RECT 1169.020 980.150 1169.620 980.290 ;
        RECT 1169.480 931.930 1169.620 980.150 ;
        RECT 1168.500 931.610 1168.760 931.930 ;
        RECT 1169.420 931.610 1169.680 931.930 ;
        RECT 1168.560 931.330 1168.700 931.610 ;
        RECT 1168.560 931.190 1169.160 931.330 ;
        RECT 1169.020 895.970 1169.160 931.190 ;
        RECT 1169.020 895.830 1169.620 895.970 ;
        RECT 1169.480 835.370 1169.620 895.830 ;
        RECT 1168.500 835.050 1168.760 835.370 ;
        RECT 1169.420 835.050 1169.680 835.370 ;
        RECT 1168.560 834.770 1168.700 835.050 ;
        RECT 1168.560 834.630 1169.160 834.770 ;
        RECT 1169.020 772.210 1169.160 834.630 ;
        RECT 1169.020 772.070 1170.080 772.210 ;
        RECT 1169.940 724.725 1170.080 772.070 ;
        RECT 1168.950 724.355 1169.230 724.725 ;
        RECT 1169.870 724.355 1170.150 724.725 ;
        RECT 1169.020 700.130 1169.160 724.355 ;
        RECT 1169.020 699.990 1169.620 700.130 ;
        RECT 1169.480 641.910 1169.620 699.990 ;
        RECT 1168.500 641.650 1168.760 641.910 ;
        RECT 1168.500 641.590 1169.160 641.650 ;
        RECT 1169.420 641.590 1169.680 641.910 ;
        RECT 1168.560 641.510 1169.160 641.590 ;
        RECT 1169.020 603.570 1169.160 641.510 ;
        RECT 1169.020 603.430 1169.620 603.570 ;
        RECT 1169.480 545.350 1169.620 603.430 ;
        RECT 1168.500 545.090 1168.760 545.350 ;
        RECT 1168.500 545.030 1169.160 545.090 ;
        RECT 1169.420 545.030 1169.680 545.350 ;
        RECT 1168.560 544.950 1169.160 545.030 ;
        RECT 1169.020 524.270 1169.160 544.950 ;
        RECT 1168.960 523.950 1169.220 524.270 ;
        RECT 1169.880 476.010 1170.140 476.330 ;
        RECT 1169.940 435.045 1170.080 476.010 ;
        RECT 1168.950 434.675 1169.230 435.045 ;
        RECT 1169.870 434.675 1170.150 435.045 ;
        RECT 1169.020 386.570 1169.160 434.675 ;
        RECT 1168.960 386.250 1169.220 386.570 ;
        RECT 1169.420 386.250 1169.680 386.570 ;
        RECT 1169.480 338.290 1169.620 386.250 ;
        RECT 1168.960 337.970 1169.220 338.290 ;
        RECT 1169.420 337.970 1169.680 338.290 ;
        RECT 1169.020 303.690 1169.160 337.970 ;
        RECT 1169.020 303.550 1169.620 303.690 ;
        RECT 1169.480 254.730 1169.620 303.550 ;
        RECT 1169.020 254.590 1169.620 254.730 ;
        RECT 1169.020 207.130 1169.160 254.590 ;
        RECT 1169.020 206.990 1169.620 207.130 ;
        RECT 1169.480 158.850 1169.620 206.990 ;
        RECT 1168.560 158.710 1169.620 158.850 ;
        RECT 1168.560 158.170 1168.700 158.710 ;
        RECT 1168.560 158.030 1169.160 158.170 ;
        RECT 1169.020 62.970 1169.160 158.030 ;
        RECT 1168.560 62.830 1169.160 62.970 ;
        RECT 1168.560 24.890 1168.700 62.830 ;
        RECT 1168.100 24.750 1168.700 24.890 ;
        RECT 1168.100 20.245 1168.240 24.750 ;
        RECT 163.390 19.875 163.670 20.245 ;
        RECT 1168.030 19.875 1168.310 20.245 ;
        RECT 163.460 2.400 163.600 19.875 ;
        RECT 163.250 -4.800 163.810 2.400 ;
      LAYER via2 ;
        RECT 1168.950 724.400 1169.230 724.680 ;
        RECT 1169.870 724.400 1170.150 724.680 ;
        RECT 1168.950 434.720 1169.230 435.000 ;
        RECT 1169.870 434.720 1170.150 435.000 ;
        RECT 163.390 19.920 163.670 20.200 ;
        RECT 1168.030 19.920 1168.310 20.200 ;
      LAYER met3 ;
        RECT 1168.925 724.690 1169.255 724.705 ;
        RECT 1169.845 724.690 1170.175 724.705 ;
        RECT 1168.925 724.390 1170.175 724.690 ;
        RECT 1168.925 724.375 1169.255 724.390 ;
        RECT 1169.845 724.375 1170.175 724.390 ;
        RECT 1168.925 435.010 1169.255 435.025 ;
        RECT 1169.845 435.010 1170.175 435.025 ;
        RECT 1168.925 434.710 1170.175 435.010 ;
        RECT 1168.925 434.695 1169.255 434.710 ;
        RECT 1169.845 434.695 1170.175 434.710 ;
        RECT 163.365 20.210 163.695 20.225 ;
        RECT 1168.005 20.210 1168.335 20.225 ;
        RECT 163.365 19.910 1168.335 20.210 ;
        RECT 163.365 19.895 163.695 19.910 ;
        RECT 1168.005 19.895 1168.335 19.910 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 196.490 1688.680 196.810 1688.740 ;
        RECT 1168.010 1688.680 1168.330 1688.740 ;
        RECT 196.490 1688.540 1168.330 1688.680 ;
        RECT 196.490 1688.480 196.810 1688.540 ;
        RECT 1168.010 1688.480 1168.330 1688.540 ;
        RECT 180.850 16.220 181.170 16.280 ;
        RECT 196.490 16.220 196.810 16.280 ;
        RECT 180.850 16.080 196.810 16.220 ;
        RECT 180.850 16.020 181.170 16.080 ;
        RECT 196.490 16.020 196.810 16.080 ;
      LAYER via ;
        RECT 196.520 1688.480 196.780 1688.740 ;
        RECT 1168.040 1688.480 1168.300 1688.740 ;
        RECT 180.880 16.020 181.140 16.280 ;
        RECT 196.520 16.020 196.780 16.280 ;
      LAYER met2 ;
        RECT 1167.940 1700.340 1168.220 1704.000 ;
        RECT 1167.940 1700.000 1168.240 1700.340 ;
        RECT 1168.100 1688.770 1168.240 1700.000 ;
        RECT 196.520 1688.450 196.780 1688.770 ;
        RECT 1168.040 1688.450 1168.300 1688.770 ;
        RECT 196.580 16.310 196.720 1688.450 ;
        RECT 180.880 15.990 181.140 16.310 ;
        RECT 196.520 15.990 196.780 16.310 ;
        RECT 180.940 2.400 181.080 15.990 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1170.310 1678.480 1170.630 1678.540 ;
        RECT 1172.150 1678.480 1172.470 1678.540 ;
        RECT 1170.310 1678.340 1172.470 1678.480 ;
        RECT 1170.310 1678.280 1170.630 1678.340 ;
        RECT 1172.150 1678.280 1172.470 1678.340 ;
        RECT 198.790 17.240 199.110 17.300 ;
        RECT 1124.770 17.240 1125.090 17.300 ;
        RECT 198.790 17.100 1125.090 17.240 ;
        RECT 198.790 17.040 199.110 17.100 ;
        RECT 1124.770 17.040 1125.090 17.100 ;
        RECT 1149.150 16.560 1149.470 16.620 ;
        RECT 1172.150 16.560 1172.470 16.620 ;
        RECT 1149.150 16.420 1172.470 16.560 ;
        RECT 1149.150 16.360 1149.470 16.420 ;
        RECT 1172.150 16.360 1172.470 16.420 ;
      LAYER via ;
        RECT 1170.340 1678.280 1170.600 1678.540 ;
        RECT 1172.180 1678.280 1172.440 1678.540 ;
        RECT 198.820 17.040 199.080 17.300 ;
        RECT 1124.800 17.040 1125.060 17.300 ;
        RECT 1149.180 16.360 1149.440 16.620 ;
        RECT 1172.180 16.360 1172.440 16.620 ;
      LAYER met2 ;
        RECT 1169.780 1700.410 1170.060 1704.000 ;
        RECT 1169.780 1700.270 1170.540 1700.410 ;
        RECT 1169.780 1700.000 1170.060 1700.270 ;
        RECT 1170.400 1678.570 1170.540 1700.270 ;
        RECT 1170.340 1678.250 1170.600 1678.570 ;
        RECT 1172.180 1678.250 1172.440 1678.570 ;
        RECT 198.820 17.010 199.080 17.330 ;
        RECT 1124.800 17.010 1125.060 17.330 ;
        RECT 198.880 2.400 199.020 17.010 ;
        RECT 1124.860 16.165 1125.000 17.010 ;
        RECT 1172.240 16.650 1172.380 1678.250 ;
        RECT 1149.180 16.330 1149.440 16.650 ;
        RECT 1172.180 16.330 1172.440 16.650 ;
        RECT 1149.240 16.165 1149.380 16.330 ;
        RECT 1124.790 15.795 1125.070 16.165 ;
        RECT 1149.170 15.795 1149.450 16.165 ;
        RECT 198.670 -4.800 199.230 2.400 ;
      LAYER via2 ;
        RECT 1124.790 15.840 1125.070 16.120 ;
        RECT 1149.170 15.840 1149.450 16.120 ;
      LAYER met3 ;
        RECT 1124.765 16.130 1125.095 16.145 ;
        RECT 1149.145 16.130 1149.475 16.145 ;
        RECT 1124.765 15.830 1149.475 16.130 ;
        RECT 1124.765 15.815 1125.095 15.830 ;
        RECT 1149.145 15.815 1149.475 15.830 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1130.825 18.105 1131.915 18.275 ;
        RECT 1130.825 17.765 1130.995 18.105 ;
        RECT 1131.745 15.215 1131.915 18.105 ;
        RECT 1131.745 15.045 1132.375 15.215 ;
      LAYER mcon ;
        RECT 1132.205 15.045 1132.375 15.215 ;
      LAYER met1 ;
        RECT 1170.310 1659.100 1170.630 1659.160 ;
        RECT 1171.690 1659.100 1172.010 1659.160 ;
        RECT 1170.310 1658.960 1172.010 1659.100 ;
        RECT 1170.310 1658.900 1170.630 1658.960 ;
        RECT 1171.690 1658.900 1172.010 1658.960 ;
        RECT 1130.765 17.920 1131.055 17.965 ;
        RECT 1125.780 17.780 1131.055 17.920 ;
        RECT 216.730 17.580 217.050 17.640 ;
        RECT 1125.780 17.580 1125.920 17.780 ;
        RECT 1130.765 17.735 1131.055 17.780 ;
        RECT 216.730 17.440 1125.920 17.580 ;
        RECT 1148.690 17.580 1149.010 17.640 ;
        RECT 1170.310 17.580 1170.630 17.640 ;
        RECT 1148.690 17.440 1170.630 17.580 ;
        RECT 216.730 17.380 217.050 17.440 ;
        RECT 1148.690 17.380 1149.010 17.440 ;
        RECT 1170.310 17.380 1170.630 17.440 ;
        RECT 1132.145 15.200 1132.435 15.245 ;
        RECT 1148.230 15.200 1148.550 15.260 ;
        RECT 1132.145 15.060 1148.550 15.200 ;
        RECT 1132.145 15.015 1132.435 15.060 ;
        RECT 1148.230 15.000 1148.550 15.060 ;
      LAYER via ;
        RECT 1170.340 1658.900 1170.600 1659.160 ;
        RECT 1171.720 1658.900 1171.980 1659.160 ;
        RECT 216.760 17.380 217.020 17.640 ;
        RECT 1148.720 17.380 1148.980 17.640 ;
        RECT 1170.340 17.380 1170.600 17.640 ;
        RECT 1148.260 15.000 1148.520 15.260 ;
      LAYER met2 ;
        RECT 1171.620 1700.340 1171.900 1704.000 ;
        RECT 1171.620 1700.000 1171.920 1700.340 ;
        RECT 1171.780 1659.190 1171.920 1700.000 ;
        RECT 1170.340 1658.870 1170.600 1659.190 ;
        RECT 1171.720 1658.870 1171.980 1659.190 ;
        RECT 1170.400 17.670 1170.540 1658.870 ;
        RECT 216.760 17.350 217.020 17.670 ;
        RECT 1148.720 17.350 1148.980 17.670 ;
        RECT 1170.340 17.350 1170.600 17.670 ;
        RECT 216.820 2.400 216.960 17.350 ;
        RECT 1148.780 16.730 1148.920 17.350 ;
        RECT 1148.320 16.590 1148.920 16.730 ;
        RECT 1148.320 15.290 1148.460 16.590 ;
        RECT 1148.260 14.970 1148.520 15.290 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1125.305 17.085 1125.475 17.935 ;
      LAYER mcon ;
        RECT 1125.305 17.765 1125.475 17.935 ;
      LAYER met1 ;
        RECT 1173.990 1658.420 1174.310 1658.480 ;
        RECT 1175.370 1658.420 1175.690 1658.480 ;
        RECT 1173.990 1658.280 1175.690 1658.420 ;
        RECT 1173.990 1658.220 1174.310 1658.280 ;
        RECT 1175.370 1658.220 1175.690 1658.280 ;
        RECT 234.670 18.260 234.990 18.320 ;
        RECT 234.670 18.120 269.400 18.260 ;
        RECT 234.670 18.060 234.990 18.120 ;
        RECT 269.260 17.920 269.400 18.120 ;
        RECT 1125.245 17.920 1125.535 17.965 ;
        RECT 269.260 17.780 1125.535 17.920 ;
        RECT 1125.245 17.735 1125.535 17.780 ;
        RECT 1125.245 17.240 1125.535 17.285 ;
        RECT 1175.370 17.240 1175.690 17.300 ;
        RECT 1125.245 17.100 1175.690 17.240 ;
        RECT 1125.245 17.055 1125.535 17.100 ;
        RECT 1175.370 17.040 1175.690 17.100 ;
      LAYER via ;
        RECT 1174.020 1658.220 1174.280 1658.480 ;
        RECT 1175.400 1658.220 1175.660 1658.480 ;
        RECT 234.700 18.060 234.960 18.320 ;
        RECT 1175.400 17.040 1175.660 17.300 ;
      LAYER met2 ;
        RECT 1173.460 1700.410 1173.740 1704.000 ;
        RECT 1173.460 1700.270 1174.220 1700.410 ;
        RECT 1173.460 1700.000 1173.740 1700.270 ;
        RECT 1174.080 1658.510 1174.220 1700.270 ;
        RECT 1174.020 1658.190 1174.280 1658.510 ;
        RECT 1175.400 1658.190 1175.660 1658.510 ;
        RECT 234.700 18.030 234.960 18.350 ;
        RECT 234.760 2.400 234.900 18.030 ;
        RECT 1175.460 17.330 1175.600 1658.190 ;
        RECT 1175.400 17.010 1175.660 17.330 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 79.190 1687.320 79.510 1687.380 ;
        RECT 1155.130 1687.320 1155.450 1687.380 ;
        RECT 79.190 1687.180 1155.450 1687.320 ;
        RECT 79.190 1687.120 79.510 1687.180 ;
        RECT 1155.130 1687.120 1155.450 1687.180 ;
        RECT 56.190 15.200 56.510 15.260 ;
        RECT 79.190 15.200 79.510 15.260 ;
        RECT 56.190 15.060 79.510 15.200 ;
        RECT 56.190 15.000 56.510 15.060 ;
        RECT 79.190 15.000 79.510 15.060 ;
      LAYER via ;
        RECT 79.220 1687.120 79.480 1687.380 ;
        RECT 1155.160 1687.120 1155.420 1687.380 ;
        RECT 56.220 15.000 56.480 15.260 ;
        RECT 79.220 15.000 79.480 15.260 ;
      LAYER met2 ;
        RECT 1155.060 1700.340 1155.340 1704.000 ;
        RECT 1155.060 1700.000 1155.360 1700.340 ;
        RECT 1155.220 1687.410 1155.360 1700.000 ;
        RECT 79.220 1687.090 79.480 1687.410 ;
        RECT 1155.160 1687.090 1155.420 1687.410 ;
        RECT 79.280 15.290 79.420 1687.090 ;
        RECT 56.220 14.970 56.480 15.290 ;
        RECT 79.220 14.970 79.480 15.290 ;
        RECT 56.280 2.400 56.420 14.970 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1157.820 1700.340 1158.100 1704.000 ;
        RECT 1157.820 1700.000 1158.120 1700.340 ;
        RECT 1157.980 18.205 1158.120 1700.000 ;
        RECT 80.130 17.835 80.410 18.205 ;
        RECT 1157.910 17.835 1158.190 18.205 ;
        RECT 80.200 2.400 80.340 17.835 ;
        RECT 79.990 -4.800 80.550 2.400 ;
      LAYER via2 ;
        RECT 80.130 17.880 80.410 18.160 ;
        RECT 1157.910 17.880 1158.190 18.160 ;
      LAYER met3 ;
        RECT 80.105 18.170 80.435 18.185 ;
        RECT 1157.885 18.170 1158.215 18.185 ;
        RECT 80.105 17.870 1158.215 18.170 ;
        RECT 80.105 17.855 80.435 17.870 ;
        RECT 1157.885 17.855 1158.215 17.870 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 141.290 1688.000 141.610 1688.060 ;
        RECT 1160.190 1688.000 1160.510 1688.060 ;
        RECT 141.290 1687.860 1160.510 1688.000 ;
        RECT 141.290 1687.800 141.610 1687.860 ;
        RECT 1160.190 1687.800 1160.510 1687.860 ;
        RECT 103.570 20.640 103.890 20.700 ;
        RECT 141.290 20.640 141.610 20.700 ;
        RECT 103.570 20.500 141.610 20.640 ;
        RECT 103.570 20.440 103.890 20.500 ;
        RECT 141.290 20.440 141.610 20.500 ;
      LAYER via ;
        RECT 141.320 1687.800 141.580 1688.060 ;
        RECT 1160.220 1687.800 1160.480 1688.060 ;
        RECT 103.600 20.440 103.860 20.700 ;
        RECT 141.320 20.440 141.580 20.700 ;
      LAYER met2 ;
        RECT 1160.120 1700.340 1160.400 1704.000 ;
        RECT 1160.120 1700.000 1160.420 1700.340 ;
        RECT 1160.280 1688.090 1160.420 1700.000 ;
        RECT 141.320 1687.770 141.580 1688.090 ;
        RECT 1160.220 1687.770 1160.480 1688.090 ;
        RECT 141.380 20.730 141.520 1687.770 ;
        RECT 103.600 20.410 103.860 20.730 ;
        RECT 141.320 20.410 141.580 20.730 ;
        RECT 103.660 2.400 103.800 20.410 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1162.490 1678.820 1162.810 1678.880 ;
        RECT 1164.790 1678.820 1165.110 1678.880 ;
        RECT 1162.490 1678.680 1165.110 1678.820 ;
        RECT 1162.490 1678.620 1162.810 1678.680 ;
        RECT 1164.790 1678.620 1165.110 1678.680 ;
      LAYER via ;
        RECT 1162.520 1678.620 1162.780 1678.880 ;
        RECT 1164.820 1678.620 1165.080 1678.880 ;
      LAYER met2 ;
        RECT 1162.420 1700.340 1162.700 1704.000 ;
        RECT 1162.420 1700.000 1162.720 1700.340 ;
        RECT 1162.580 1678.910 1162.720 1700.000 ;
        RECT 1162.520 1678.590 1162.780 1678.910 ;
        RECT 1164.820 1678.590 1165.080 1678.910 ;
        RECT 1164.880 19.565 1165.020 1678.590 ;
        RECT 127.510 19.195 127.790 19.565 ;
        RECT 1164.810 19.195 1165.090 19.565 ;
        RECT 127.580 2.400 127.720 19.195 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 127.510 19.240 127.790 19.520 ;
        RECT 1164.810 19.240 1165.090 19.520 ;
      LAYER met3 ;
        RECT 127.485 19.530 127.815 19.545 ;
        RECT 1164.785 19.530 1165.115 19.545 ;
        RECT 127.485 19.230 1165.115 19.530 ;
        RECT 127.485 19.215 127.815 19.230 ;
        RECT 1164.785 19.215 1165.115 19.230 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 51.590 1686.980 51.910 1687.040 ;
        RECT 1152.370 1686.980 1152.690 1687.040 ;
        RECT 51.590 1686.840 1152.690 1686.980 ;
        RECT 51.590 1686.780 51.910 1686.840 ;
        RECT 1152.370 1686.780 1152.690 1686.840 ;
        RECT 26.290 17.240 26.610 17.300 ;
        RECT 51.590 17.240 51.910 17.300 ;
        RECT 26.290 17.100 51.910 17.240 ;
        RECT 26.290 17.040 26.610 17.100 ;
        RECT 51.590 17.040 51.910 17.100 ;
      LAYER via ;
        RECT 51.620 1686.780 51.880 1687.040 ;
        RECT 1152.400 1686.780 1152.660 1687.040 ;
        RECT 26.320 17.040 26.580 17.300 ;
        RECT 51.620 17.040 51.880 17.300 ;
      LAYER met2 ;
        RECT 1152.300 1700.340 1152.580 1704.000 ;
        RECT 1152.300 1700.000 1152.600 1700.340 ;
        RECT 1152.460 1687.070 1152.600 1700.000 ;
        RECT 51.620 1686.750 51.880 1687.070 ;
        RECT 1152.400 1686.750 1152.660 1687.070 ;
        RECT 51.680 17.330 51.820 1686.750 ;
        RECT 26.320 17.010 26.580 17.330 ;
        RECT 51.620 17.010 51.880 17.330 ;
        RECT 26.380 2.400 26.520 17.010 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1152.830 1677.460 1153.150 1677.520 ;
        RECT 1155.590 1677.460 1155.910 1677.520 ;
        RECT 1152.830 1677.320 1155.910 1677.460 ;
        RECT 1152.830 1677.260 1153.150 1677.320 ;
        RECT 1155.590 1677.260 1155.910 1677.320 ;
      LAYER via ;
        RECT 1152.860 1677.260 1153.120 1677.520 ;
        RECT 1155.620 1677.260 1155.880 1677.520 ;
      LAYER met2 ;
        RECT 1152.760 1700.340 1153.040 1704.000 ;
        RECT 1152.760 1700.000 1153.060 1700.340 ;
        RECT 1152.920 1677.550 1153.060 1700.000 ;
        RECT 1152.860 1677.230 1153.120 1677.550 ;
        RECT 1155.620 1677.230 1155.880 1677.550 ;
        RECT 1155.680 16.845 1155.820 1677.230 ;
        RECT 32.290 16.475 32.570 16.845 ;
        RECT 1155.610 16.475 1155.890 16.845 ;
        RECT 32.360 2.400 32.500 16.475 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 32.290 16.520 32.570 16.800 ;
        RECT 1155.610 16.520 1155.890 16.800 ;
      LAYER met3 ;
        RECT 32.265 16.810 32.595 16.825 ;
        RECT 1155.585 16.810 1155.915 16.825 ;
        RECT 32.265 16.510 1155.915 16.810 ;
        RECT 32.265 16.495 32.595 16.510 ;
        RECT 1155.585 16.495 1155.915 16.510 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 -9.220 367.020 3528.900 ;
        RECT 544.020 -9.220 547.020 3528.900 ;
        RECT 724.020 -9.220 727.020 3528.900 ;
        RECT 904.020 -9.220 907.020 3528.900 ;
        RECT 1084.020 -9.220 1087.020 3528.900 ;
        RECT 1264.020 -9.220 1267.020 3528.900 ;
        RECT 1444.020 -9.220 1447.020 3528.900 ;
        RECT 1624.020 -9.220 1627.020 3528.900 ;
        RECT 1804.020 -9.220 1807.020 3528.900 ;
        RECT 1984.020 -9.220 1987.020 3528.900 ;
        RECT 2164.020 -9.220 2167.020 3528.900 ;
        RECT 2344.020 -9.220 2347.020 3528.900 ;
        RECT 2524.020 -9.220 2527.020 3528.900 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 -9.220 457.020 3528.900 ;
        RECT 634.020 -9.220 637.020 3528.900 ;
        RECT 814.020 -9.220 817.020 3528.900 ;
        RECT 994.020 -9.220 997.020 3528.900 ;
        RECT 1174.020 -9.220 1177.020 3528.900 ;
        RECT 1354.020 -9.220 1357.020 3528.900 ;
        RECT 1534.020 -9.220 1537.020 3528.900 ;
        RECT 1714.020 -9.220 1717.020 3528.900 ;
        RECT 1894.020 -9.220 1897.020 3528.900 ;
        RECT 2074.020 -9.220 2077.020 3528.900 ;
        RECT 2254.020 -9.220 2257.020 3528.900 ;
        RECT 2434.020 -9.220 2437.020 3528.900 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 -18.420 385.020 3538.100 ;
        RECT 562.020 -18.420 565.020 3538.100 ;
        RECT 742.020 -18.420 745.020 3538.100 ;
        RECT 922.020 -18.420 925.020 3538.100 ;
        RECT 1102.020 -18.420 1105.020 3538.100 ;
        RECT 1282.020 -18.420 1285.020 3538.100 ;
        RECT 1462.020 -18.420 1465.020 3538.100 ;
        RECT 1642.020 -18.420 1645.020 3538.100 ;
        RECT 1822.020 -18.420 1825.020 3538.100 ;
        RECT 2002.020 -18.420 2005.020 3538.100 ;
        RECT 2182.020 -18.420 2185.020 3538.100 ;
        RECT 2362.020 -18.420 2365.020 3538.100 ;
        RECT 2542.020 -18.420 2545.020 3538.100 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1102.930 2009.090 1104.110 2010.270 ;
        RECT 1102.930 2007.490 1104.110 2008.670 ;
        RECT 1102.930 1829.090 1104.110 1830.270 ;
        RECT 1102.930 1827.490 1104.110 1828.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1282.930 2009.090 1284.110 2010.270 ;
        RECT 1282.930 2007.490 1284.110 2008.670 ;
        RECT 1282.930 1829.090 1284.110 1830.270 ;
        RECT 1282.930 1827.490 1284.110 1828.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1102.020 2010.380 1105.020 2010.390 ;
        RECT 1282.020 2010.380 1285.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1102.020 2007.370 1105.020 2007.380 ;
        RECT 1282.020 2007.370 1285.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1102.020 1830.380 1105.020 1830.390 ;
        RECT 1282.020 1830.380 1285.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1102.020 1827.370 1105.020 1827.380 ;
        RECT 1282.020 1827.370 1285.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 -18.420 475.020 3538.100 ;
        RECT 652.020 -18.420 655.020 3538.100 ;
        RECT 832.020 -18.420 835.020 3538.100 ;
        RECT 1012.020 -18.420 1015.020 3538.100 ;
        RECT 1192.020 -18.420 1195.020 3538.100 ;
        RECT 1372.020 -18.420 1375.020 3538.100 ;
        RECT 1552.020 -18.420 1555.020 3538.100 ;
        RECT 1732.020 -18.420 1735.020 3538.100 ;
        RECT 1912.020 -18.420 1915.020 3538.100 ;
        RECT 2092.020 -18.420 2095.020 3538.100 ;
        RECT 2272.020 -18.420 2275.020 3538.100 ;
        RECT 2452.020 -18.420 2455.020 3538.100 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1012.930 1919.090 1014.110 1920.270 ;
        RECT 1012.930 1917.490 1014.110 1918.670 ;
        RECT 1012.930 1739.090 1014.110 1740.270 ;
        RECT 1012.930 1737.490 1014.110 1738.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1192.930 1919.090 1194.110 1920.270 ;
        RECT 1192.930 1917.490 1194.110 1918.670 ;
        RECT 1192.930 1739.090 1194.110 1740.270 ;
        RECT 1192.930 1737.490 1194.110 1738.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1012.020 1920.380 1015.020 1920.390 ;
        RECT 1192.020 1920.380 1195.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1012.020 1917.370 1015.020 1917.380 ;
        RECT 1192.020 1917.370 1195.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1012.020 1740.380 1015.020 1740.390 ;
        RECT 1192.020 1740.380 1195.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1012.020 1737.370 1015.020 1737.380 ;
        RECT 1192.020 1737.370 1195.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 -27.620 403.020 3547.300 ;
        RECT 580.020 -27.620 583.020 3547.300 ;
        RECT 760.020 -27.620 763.020 3547.300 ;
        RECT 940.020 -27.620 943.020 3547.300 ;
        RECT 1120.020 -27.620 1123.020 3547.300 ;
        RECT 1300.020 -27.620 1303.020 3547.300 ;
        RECT 1480.020 -27.620 1483.020 3547.300 ;
        RECT 1660.020 -27.620 1663.020 3547.300 ;
        RECT 1840.020 -27.620 1843.020 3547.300 ;
        RECT 2020.020 -27.620 2023.020 3547.300 ;
        RECT 2200.020 -27.620 2203.020 3547.300 ;
        RECT 2380.020 -27.620 2383.020 3547.300 ;
        RECT 2560.020 -27.620 2563.020 3547.300 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1120.930 2027.090 1122.110 2028.270 ;
        RECT 1120.930 2025.490 1122.110 2026.670 ;
        RECT 1120.930 1847.090 1122.110 1848.270 ;
        RECT 1120.930 1845.490 1122.110 1846.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1300.930 2027.090 1302.110 2028.270 ;
        RECT 1300.930 2025.490 1302.110 2026.670 ;
        RECT 1300.930 1847.090 1302.110 1848.270 ;
        RECT 1300.930 1845.490 1302.110 1846.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1120.020 2028.380 1123.020 2028.390 ;
        RECT 1300.020 2028.380 1303.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1120.020 2025.370 1123.020 2025.380 ;
        RECT 1300.020 2025.370 1303.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1120.020 1848.380 1123.020 1848.390 ;
        RECT 1300.020 1848.380 1303.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1120.020 1845.370 1123.020 1845.380 ;
        RECT 1300.020 1845.370 1303.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 -27.620 313.020 3547.300 ;
        RECT 490.020 -27.620 493.020 3547.300 ;
        RECT 670.020 -27.620 673.020 3547.300 ;
        RECT 850.020 -27.620 853.020 3547.300 ;
        RECT 1030.020 -27.620 1033.020 3547.300 ;
        RECT 1210.020 -27.620 1213.020 3547.300 ;
        RECT 1390.020 -27.620 1393.020 3547.300 ;
        RECT 1570.020 -27.620 1573.020 3547.300 ;
        RECT 1750.020 -27.620 1753.020 3547.300 ;
        RECT 1930.020 -27.620 1933.020 3547.300 ;
        RECT 2110.020 -27.620 2113.020 3547.300 ;
        RECT 2290.020 -27.620 2293.020 3547.300 ;
        RECT 2470.020 -27.620 2473.020 3547.300 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1030.930 2657.090 1032.110 2658.270 ;
        RECT 1030.930 2655.490 1032.110 2656.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1030.930 1937.090 1032.110 1938.270 ;
        RECT 1030.930 1935.490 1032.110 1936.670 ;
        RECT 1030.930 1757.090 1032.110 1758.270 ;
        RECT 1030.930 1755.490 1032.110 1756.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1210.930 1937.090 1212.110 1938.270 ;
        RECT 1210.930 1935.490 1212.110 1936.670 ;
        RECT 1210.930 1757.090 1212.110 1758.270 ;
        RECT 1210.930 1755.490 1212.110 1756.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1570.930 2837.090 1572.110 2838.270 ;
        RECT 1570.930 2835.490 1572.110 2836.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1750.930 2837.090 1752.110 2838.270 ;
        RECT 1750.930 2835.490 1752.110 2836.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 1930.930 1757.090 1932.110 1758.270 ;
        RECT 1930.930 1755.490 1932.110 1756.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1570.020 2838.380 1573.020 2838.390 ;
        RECT 1750.020 2838.380 1753.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1570.020 2835.370 1573.020 2835.380 ;
        RECT 1750.020 2835.370 1753.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1030.020 2658.380 1033.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1030.020 2655.370 1033.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1030.020 1938.380 1033.020 1938.390 ;
        RECT 1210.020 1938.380 1213.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1030.020 1935.370 1033.020 1935.380 ;
        RECT 1210.020 1935.370 1213.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1030.020 1758.380 1033.020 1758.390 ;
        RECT 1210.020 1758.380 1213.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 1930.020 1758.380 1933.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1030.020 1755.370 1033.020 1755.380 ;
        RECT 1210.020 1755.370 1213.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 1930.020 1755.370 1933.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 -36.820 421.020 3556.500 ;
        RECT 598.020 -36.820 601.020 3556.500 ;
        RECT 778.020 -36.820 781.020 3556.500 ;
        RECT 958.020 -36.820 961.020 3556.500 ;
        RECT 1138.020 -36.820 1141.020 3556.500 ;
        RECT 1318.020 -36.820 1321.020 3556.500 ;
        RECT 1498.020 -36.820 1501.020 3556.500 ;
        RECT 1678.020 -36.820 1681.020 3556.500 ;
        RECT 1858.020 -36.820 1861.020 3556.500 ;
        RECT 2038.020 -36.820 2041.020 3556.500 ;
        RECT 2218.020 -36.820 2221.020 3556.500 ;
        RECT 2398.020 -36.820 2401.020 3556.500 ;
        RECT 2578.020 -36.820 2581.020 3556.500 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1138.930 2045.090 1140.110 2046.270 ;
        RECT 1138.930 2043.490 1140.110 2044.670 ;
        RECT 1138.930 1865.090 1140.110 1866.270 ;
        RECT 1138.930 1863.490 1140.110 1864.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1318.930 2045.090 1320.110 2046.270 ;
        RECT 1318.930 2043.490 1320.110 2044.670 ;
        RECT 1318.930 1865.090 1320.110 1866.270 ;
        RECT 1318.930 1863.490 1320.110 1864.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1138.020 2046.380 1141.020 2046.390 ;
        RECT 1318.020 2046.380 1321.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1138.020 2043.370 1141.020 2043.380 ;
        RECT 1318.020 2043.370 1321.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1138.020 1866.380 1141.020 1866.390 ;
        RECT 1318.020 1866.380 1321.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1138.020 1863.370 1141.020 1863.380 ;
        RECT 1318.020 1863.370 1321.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 -36.820 331.020 3556.500 ;
        RECT 508.020 -36.820 511.020 3556.500 ;
        RECT 688.020 -36.820 691.020 3556.500 ;
        RECT 868.020 -36.820 871.020 3556.500 ;
        RECT 1048.020 -36.820 1051.020 3556.500 ;
        RECT 1228.020 -36.820 1231.020 3556.500 ;
        RECT 1408.020 -36.820 1411.020 3556.500 ;
        RECT 1588.020 -36.820 1591.020 3556.500 ;
        RECT 1768.020 -36.820 1771.020 3556.500 ;
        RECT 1948.020 -36.820 1951.020 3556.500 ;
        RECT 2128.020 -36.820 2131.020 3556.500 ;
        RECT 2308.020 -36.820 2311.020 3556.500 ;
        RECT 2488.020 -36.820 2491.020 3556.500 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1048.930 2675.090 1050.110 2676.270 ;
        RECT 1048.930 2673.490 1050.110 2674.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1048.930 1955.090 1050.110 1956.270 ;
        RECT 1048.930 1953.490 1050.110 1954.670 ;
        RECT 1048.930 1775.090 1050.110 1776.270 ;
        RECT 1048.930 1773.490 1050.110 1774.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1228.930 1955.090 1230.110 1956.270 ;
        RECT 1228.930 1953.490 1230.110 1954.670 ;
        RECT 1228.930 1775.090 1230.110 1776.270 ;
        RECT 1228.930 1773.490 1230.110 1774.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1588.930 2855.090 1590.110 2856.270 ;
        RECT 1588.930 2853.490 1590.110 2854.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1768.930 2855.090 1770.110 2856.270 ;
        RECT 1768.930 2853.490 1770.110 2854.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 1948.930 1775.090 1950.110 1776.270 ;
        RECT 1948.930 1773.490 1950.110 1774.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1588.020 2856.380 1591.020 2856.390 ;
        RECT 1768.020 2856.380 1771.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1588.020 2853.370 1591.020 2853.380 ;
        RECT 1768.020 2853.370 1771.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1048.020 2676.380 1051.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1048.020 2673.370 1051.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1048.020 1956.380 1051.020 1956.390 ;
        RECT 1228.020 1956.380 1231.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1048.020 1953.370 1051.020 1953.380 ;
        RECT 1228.020 1953.370 1231.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1048.020 1776.380 1051.020 1776.390 ;
        RECT 1228.020 1776.380 1231.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 1948.020 1776.380 1951.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1048.020 1773.370 1051.020 1773.380 ;
        RECT 1228.020 1773.370 1231.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 1948.020 1773.370 1951.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 1155.430 1710.795 1444.310 1988.405 ;
      LAYER met1 ;
        RECT 1150.900 1704.460 1448.840 1989.980 ;
      LAYER met2 ;
        RECT 1151.480 1995.720 1152.940 1996.000 ;
        RECT 1153.780 1995.720 1155.700 1996.000 ;
        RECT 1156.540 1995.720 1158.460 1996.000 ;
        RECT 1159.300 1995.720 1160.760 1996.000 ;
        RECT 1161.600 1995.720 1163.520 1996.000 ;
        RECT 1164.360 1995.720 1166.280 1996.000 ;
        RECT 1167.120 1995.720 1169.040 1996.000 ;
        RECT 1169.880 1995.720 1171.340 1996.000 ;
        RECT 1172.180 1995.720 1174.100 1996.000 ;
        RECT 1174.940 1995.720 1176.860 1996.000 ;
        RECT 1177.700 1995.720 1179.160 1996.000 ;
        RECT 1180.000 1995.720 1181.920 1996.000 ;
        RECT 1182.760 1995.720 1184.680 1996.000 ;
        RECT 1185.520 1995.720 1187.440 1996.000 ;
        RECT 1188.280 1995.720 1189.740 1996.000 ;
        RECT 1190.580 1995.720 1192.500 1996.000 ;
        RECT 1193.340 1995.720 1195.260 1996.000 ;
        RECT 1196.100 1995.720 1197.560 1996.000 ;
        RECT 1198.400 1995.720 1200.320 1996.000 ;
        RECT 1201.160 1995.720 1203.080 1996.000 ;
        RECT 1203.920 1995.720 1205.840 1996.000 ;
        RECT 1206.680 1995.720 1208.140 1996.000 ;
        RECT 1208.980 1995.720 1210.900 1996.000 ;
        RECT 1211.740 1995.720 1213.660 1996.000 ;
        RECT 1214.500 1995.720 1215.960 1996.000 ;
        RECT 1216.800 1995.720 1218.720 1996.000 ;
        RECT 1219.560 1995.720 1221.480 1996.000 ;
        RECT 1222.320 1995.720 1224.240 1996.000 ;
        RECT 1225.080 1995.720 1226.540 1996.000 ;
        RECT 1227.380 1995.720 1229.300 1996.000 ;
        RECT 1230.140 1995.720 1232.060 1996.000 ;
        RECT 1232.900 1995.720 1234.820 1996.000 ;
        RECT 1235.660 1995.720 1237.120 1996.000 ;
        RECT 1237.960 1995.720 1239.880 1996.000 ;
        RECT 1240.720 1995.720 1242.640 1996.000 ;
        RECT 1243.480 1995.720 1244.940 1996.000 ;
        RECT 1245.780 1995.720 1247.700 1996.000 ;
        RECT 1248.540 1995.720 1250.460 1996.000 ;
        RECT 1251.300 1995.720 1253.220 1996.000 ;
        RECT 1254.060 1995.720 1255.520 1996.000 ;
        RECT 1256.360 1995.720 1258.280 1996.000 ;
        RECT 1259.120 1995.720 1261.040 1996.000 ;
        RECT 1261.880 1995.720 1263.340 1996.000 ;
        RECT 1264.180 1995.720 1266.100 1996.000 ;
        RECT 1266.940 1995.720 1268.860 1996.000 ;
        RECT 1269.700 1995.720 1271.620 1996.000 ;
        RECT 1272.460 1995.720 1273.920 1996.000 ;
        RECT 1274.760 1995.720 1276.680 1996.000 ;
        RECT 1277.520 1995.720 1279.440 1996.000 ;
        RECT 1280.280 1995.720 1281.740 1996.000 ;
        RECT 1282.580 1995.720 1284.500 1996.000 ;
        RECT 1285.340 1995.720 1287.260 1996.000 ;
        RECT 1288.100 1995.720 1290.020 1996.000 ;
        RECT 1290.860 1995.720 1292.320 1996.000 ;
        RECT 1293.160 1995.720 1295.080 1996.000 ;
        RECT 1295.920 1995.720 1297.840 1996.000 ;
        RECT 1298.680 1995.720 1300.600 1996.000 ;
        RECT 1301.440 1995.720 1302.900 1996.000 ;
        RECT 1303.740 1995.720 1305.660 1996.000 ;
        RECT 1306.500 1995.720 1308.420 1996.000 ;
        RECT 1309.260 1995.720 1310.720 1996.000 ;
        RECT 1311.560 1995.720 1313.480 1996.000 ;
        RECT 1314.320 1995.720 1316.240 1996.000 ;
        RECT 1317.080 1995.720 1319.000 1996.000 ;
        RECT 1319.840 1995.720 1321.300 1996.000 ;
        RECT 1322.140 1995.720 1324.060 1996.000 ;
        RECT 1324.900 1995.720 1326.820 1996.000 ;
        RECT 1327.660 1995.720 1329.120 1996.000 ;
        RECT 1329.960 1995.720 1331.880 1996.000 ;
        RECT 1332.720 1995.720 1334.640 1996.000 ;
        RECT 1335.480 1995.720 1337.400 1996.000 ;
        RECT 1338.240 1995.720 1339.700 1996.000 ;
        RECT 1340.540 1995.720 1342.460 1996.000 ;
        RECT 1343.300 1995.720 1345.220 1996.000 ;
        RECT 1346.060 1995.720 1347.520 1996.000 ;
        RECT 1348.360 1995.720 1350.280 1996.000 ;
        RECT 1351.120 1995.720 1353.040 1996.000 ;
        RECT 1353.880 1995.720 1355.800 1996.000 ;
        RECT 1356.640 1995.720 1358.100 1996.000 ;
        RECT 1358.940 1995.720 1360.860 1996.000 ;
        RECT 1361.700 1995.720 1363.620 1996.000 ;
        RECT 1364.460 1995.720 1365.920 1996.000 ;
        RECT 1366.760 1995.720 1368.680 1996.000 ;
        RECT 1369.520 1995.720 1371.440 1996.000 ;
        RECT 1372.280 1995.720 1374.200 1996.000 ;
        RECT 1375.040 1995.720 1376.500 1996.000 ;
        RECT 1377.340 1995.720 1379.260 1996.000 ;
        RECT 1380.100 1995.720 1382.020 1996.000 ;
        RECT 1382.860 1995.720 1384.780 1996.000 ;
        RECT 1385.620 1995.720 1387.080 1996.000 ;
        RECT 1387.920 1995.720 1389.840 1996.000 ;
        RECT 1390.680 1995.720 1392.600 1996.000 ;
        RECT 1393.440 1995.720 1394.900 1996.000 ;
        RECT 1395.740 1995.720 1397.660 1996.000 ;
        RECT 1398.500 1995.720 1400.420 1996.000 ;
        RECT 1401.260 1995.720 1403.180 1996.000 ;
        RECT 1404.020 1995.720 1405.480 1996.000 ;
        RECT 1406.320 1995.720 1408.240 1996.000 ;
        RECT 1409.080 1995.720 1411.000 1996.000 ;
        RECT 1411.840 1995.720 1413.300 1996.000 ;
        RECT 1414.140 1995.720 1416.060 1996.000 ;
        RECT 1416.900 1995.720 1418.820 1996.000 ;
        RECT 1419.660 1995.720 1421.580 1996.000 ;
        RECT 1422.420 1995.720 1423.880 1996.000 ;
        RECT 1424.720 1995.720 1426.640 1996.000 ;
        RECT 1427.480 1995.720 1429.400 1996.000 ;
        RECT 1430.240 1995.720 1431.700 1996.000 ;
        RECT 1432.540 1995.720 1434.460 1996.000 ;
        RECT 1435.300 1995.720 1437.220 1996.000 ;
        RECT 1438.060 1995.720 1439.980 1996.000 ;
        RECT 1440.820 1995.720 1442.280 1996.000 ;
        RECT 1443.120 1995.720 1445.040 1996.000 ;
        RECT 1445.880 1995.720 1447.800 1996.000 ;
        RECT 1448.640 1995.720 1448.810 1996.000 ;
        RECT 1150.930 1704.280 1448.810 1995.720 ;
        RECT 1151.940 1704.000 1152.020 1704.280 ;
        RECT 1153.780 1704.000 1153.860 1704.280 ;
        RECT 1155.620 1704.000 1155.700 1704.280 ;
        RECT 1157.460 1704.000 1157.540 1704.280 ;
        RECT 1159.300 1704.000 1159.380 1704.280 ;
        RECT 1161.140 1704.000 1161.220 1704.280 ;
        RECT 1162.980 1704.000 1163.060 1704.280 ;
        RECT 1164.820 1704.000 1164.900 1704.280 ;
        RECT 1166.660 1704.000 1166.740 1704.280 ;
        RECT 1168.500 1704.000 1168.580 1704.280 ;
        RECT 1170.340 1704.000 1170.420 1704.280 ;
        RECT 1172.180 1704.000 1172.260 1704.280 ;
        RECT 1174.020 1704.000 1174.100 1704.280 ;
        RECT 1175.860 1704.000 1175.940 1704.280 ;
        RECT 1177.700 1704.000 1177.780 1704.280 ;
        RECT 1179.540 1704.000 1179.620 1704.280 ;
        RECT 1181.380 1704.000 1181.460 1704.280 ;
        RECT 1183.220 1704.000 1183.300 1704.280 ;
        RECT 1185.060 1704.000 1185.140 1704.280 ;
        RECT 1186.900 1704.000 1186.980 1704.280 ;
        RECT 1188.740 1704.000 1188.820 1704.280 ;
        RECT 1190.580 1704.000 1190.660 1704.280 ;
        RECT 1192.420 1704.000 1192.500 1704.280 ;
        RECT 1194.260 1704.000 1194.340 1704.280 ;
        RECT 1196.100 1704.000 1196.180 1704.280 ;
        RECT 1197.940 1704.000 1198.020 1704.280 ;
        RECT 1199.780 1704.000 1199.860 1704.280 ;
        RECT 1201.620 1704.000 1201.700 1704.280 ;
        RECT 1203.460 1704.000 1203.540 1704.280 ;
        RECT 1205.300 1704.000 1205.380 1704.280 ;
        RECT 1207.140 1704.000 1207.220 1704.280 ;
        RECT 1208.980 1704.000 1209.060 1704.280 ;
        RECT 1210.820 1704.000 1210.900 1704.280 ;
        RECT 1212.660 1704.000 1212.740 1704.280 ;
        RECT 1214.500 1704.000 1214.580 1704.280 ;
        RECT 1216.340 1704.000 1216.420 1704.280 ;
        RECT 1218.180 1704.000 1218.260 1704.280 ;
        RECT 1220.020 1704.000 1220.100 1704.280 ;
        RECT 1221.860 1704.000 1221.940 1704.280 ;
        RECT 1223.700 1704.000 1223.780 1704.280 ;
        RECT 1226.000 1704.000 1226.080 1704.280 ;
        RECT 1227.840 1704.000 1227.920 1704.280 ;
        RECT 1229.680 1704.000 1229.760 1704.280 ;
        RECT 1231.520 1704.000 1231.600 1704.280 ;
        RECT 1233.360 1704.000 1233.440 1704.280 ;
        RECT 1235.200 1704.000 1235.280 1704.280 ;
        RECT 1237.040 1704.000 1237.120 1704.280 ;
        RECT 1238.880 1704.000 1238.960 1704.280 ;
        RECT 1240.720 1704.000 1240.800 1704.280 ;
        RECT 1242.560 1704.000 1242.640 1704.280 ;
        RECT 1244.400 1704.000 1244.480 1704.280 ;
        RECT 1246.240 1704.000 1246.320 1704.280 ;
        RECT 1248.080 1704.000 1248.160 1704.280 ;
        RECT 1249.920 1704.000 1250.000 1704.280 ;
        RECT 1251.760 1704.000 1251.840 1704.280 ;
        RECT 1253.600 1704.000 1253.680 1704.280 ;
        RECT 1255.440 1704.000 1255.520 1704.280 ;
        RECT 1257.280 1704.000 1257.360 1704.280 ;
        RECT 1259.120 1704.000 1259.200 1704.280 ;
        RECT 1260.960 1704.000 1261.040 1704.280 ;
        RECT 1262.800 1704.000 1262.880 1704.280 ;
        RECT 1264.640 1704.000 1264.720 1704.280 ;
        RECT 1266.480 1704.000 1266.560 1704.280 ;
        RECT 1268.320 1704.000 1268.400 1704.280 ;
        RECT 1270.160 1704.000 1270.240 1704.280 ;
        RECT 1272.000 1704.000 1272.080 1704.280 ;
        RECT 1273.840 1704.000 1273.920 1704.280 ;
        RECT 1275.680 1704.000 1275.760 1704.280 ;
        RECT 1277.520 1704.000 1277.600 1704.280 ;
        RECT 1279.360 1704.000 1279.440 1704.280 ;
        RECT 1281.200 1704.000 1281.280 1704.280 ;
        RECT 1283.040 1704.000 1283.120 1704.280 ;
        RECT 1284.880 1704.000 1284.960 1704.280 ;
        RECT 1286.720 1704.000 1286.800 1704.280 ;
        RECT 1288.560 1704.000 1288.640 1704.280 ;
        RECT 1290.400 1704.000 1290.480 1704.280 ;
        RECT 1292.240 1704.000 1292.320 1704.280 ;
        RECT 1294.080 1704.000 1294.160 1704.280 ;
        RECT 1295.920 1704.000 1296.000 1704.280 ;
        RECT 1297.760 1704.000 1297.840 1704.280 ;
        RECT 1299.600 1704.000 1299.680 1704.280 ;
        RECT 1301.900 1704.000 1301.980 1704.280 ;
        RECT 1303.740 1704.000 1303.820 1704.280 ;
        RECT 1305.580 1704.000 1305.660 1704.280 ;
        RECT 1307.420 1704.000 1307.500 1704.280 ;
        RECT 1309.260 1704.000 1309.340 1704.280 ;
        RECT 1311.100 1704.000 1311.180 1704.280 ;
        RECT 1312.940 1704.000 1313.020 1704.280 ;
        RECT 1314.780 1704.000 1314.860 1704.280 ;
        RECT 1316.620 1704.000 1316.700 1704.280 ;
        RECT 1318.460 1704.000 1318.540 1704.280 ;
        RECT 1320.300 1704.000 1320.380 1704.280 ;
        RECT 1322.140 1704.000 1322.220 1704.280 ;
        RECT 1323.980 1704.000 1324.060 1704.280 ;
        RECT 1325.820 1704.000 1325.900 1704.280 ;
        RECT 1327.660 1704.000 1327.740 1704.280 ;
        RECT 1329.500 1704.000 1329.580 1704.280 ;
        RECT 1331.340 1704.000 1331.420 1704.280 ;
        RECT 1333.180 1704.000 1333.260 1704.280 ;
        RECT 1335.020 1704.000 1335.100 1704.280 ;
        RECT 1336.860 1704.000 1336.940 1704.280 ;
        RECT 1338.700 1704.000 1338.780 1704.280 ;
        RECT 1340.540 1704.000 1340.620 1704.280 ;
        RECT 1342.380 1704.000 1342.460 1704.280 ;
        RECT 1344.220 1704.000 1344.300 1704.280 ;
        RECT 1346.060 1704.000 1346.140 1704.280 ;
        RECT 1347.900 1704.000 1347.980 1704.280 ;
        RECT 1349.740 1704.000 1349.820 1704.280 ;
        RECT 1351.580 1704.000 1351.660 1704.280 ;
        RECT 1353.420 1704.000 1353.500 1704.280 ;
        RECT 1355.260 1704.000 1355.340 1704.280 ;
        RECT 1357.100 1704.000 1357.180 1704.280 ;
        RECT 1358.940 1704.000 1359.020 1704.280 ;
        RECT 1360.780 1704.000 1360.860 1704.280 ;
        RECT 1362.620 1704.000 1362.700 1704.280 ;
        RECT 1364.460 1704.000 1364.540 1704.280 ;
        RECT 1366.300 1704.000 1366.380 1704.280 ;
        RECT 1368.140 1704.000 1368.220 1704.280 ;
        RECT 1369.980 1704.000 1370.060 1704.280 ;
        RECT 1371.820 1704.000 1371.900 1704.280 ;
        RECT 1373.660 1704.000 1373.740 1704.280 ;
        RECT 1375.960 1704.000 1376.040 1704.280 ;
        RECT 1377.800 1704.000 1377.880 1704.280 ;
        RECT 1379.640 1704.000 1379.720 1704.280 ;
        RECT 1381.480 1704.000 1381.560 1704.280 ;
        RECT 1383.320 1704.000 1383.400 1704.280 ;
        RECT 1385.160 1704.000 1385.240 1704.280 ;
        RECT 1387.000 1704.000 1387.080 1704.280 ;
        RECT 1388.840 1704.000 1388.920 1704.280 ;
        RECT 1390.680 1704.000 1390.760 1704.280 ;
        RECT 1392.520 1704.000 1392.600 1704.280 ;
        RECT 1394.360 1704.000 1394.440 1704.280 ;
        RECT 1396.200 1704.000 1396.280 1704.280 ;
        RECT 1398.040 1704.000 1398.120 1704.280 ;
        RECT 1399.880 1704.000 1399.960 1704.280 ;
        RECT 1401.720 1704.000 1401.800 1704.280 ;
        RECT 1403.560 1704.000 1403.640 1704.280 ;
        RECT 1405.400 1704.000 1405.480 1704.280 ;
        RECT 1407.240 1704.000 1407.320 1704.280 ;
        RECT 1409.080 1704.000 1409.160 1704.280 ;
        RECT 1410.920 1704.000 1411.000 1704.280 ;
        RECT 1412.760 1704.000 1412.840 1704.280 ;
        RECT 1414.600 1704.000 1414.680 1704.280 ;
        RECT 1416.440 1704.000 1416.520 1704.280 ;
        RECT 1418.280 1704.000 1418.360 1704.280 ;
        RECT 1420.120 1704.000 1420.200 1704.280 ;
        RECT 1421.960 1704.000 1422.040 1704.280 ;
        RECT 1423.800 1704.000 1423.880 1704.280 ;
        RECT 1425.640 1704.000 1425.720 1704.280 ;
        RECT 1427.480 1704.000 1427.560 1704.280 ;
        RECT 1429.320 1704.000 1429.400 1704.280 ;
        RECT 1431.160 1704.000 1431.240 1704.280 ;
        RECT 1433.000 1704.000 1433.080 1704.280 ;
        RECT 1434.840 1704.000 1434.920 1704.280 ;
        RECT 1436.680 1704.000 1436.760 1704.280 ;
        RECT 1438.520 1704.000 1438.600 1704.280 ;
        RECT 1440.360 1704.000 1440.440 1704.280 ;
        RECT 1442.200 1704.000 1442.280 1704.280 ;
        RECT 1444.040 1704.000 1444.120 1704.280 ;
        RECT 1445.880 1704.000 1445.960 1704.280 ;
        RECT 1447.720 1704.000 1447.800 1704.280 ;
      LAYER met3 ;
        RECT 1154.575 1704.255 1434.585 1988.485 ;
      LAYER met4 ;
        RECT 1170.950 1710.640 1172.550 1988.560 ;
      LAYER met4 ;
        RECT 1196.205 1710.640 1210.020 1988.560 ;
        RECT 1213.020 1710.640 1228.020 1988.560 ;
        RECT 1231.020 1710.640 1247.350 1988.560 ;
      LAYER met4 ;
        RECT 1247.750 1710.640 1249.350 1988.560 ;
      LAYER met4 ;
        RECT 1249.750 1710.640 1264.020 1988.560 ;
        RECT 1267.020 1710.640 1282.020 1988.560 ;
        RECT 1285.020 1710.640 1300.020 1988.560 ;
        RECT 1303.020 1710.640 1318.020 1988.560 ;
        RECT 1321.020 1710.640 1354.020 1988.560 ;
        RECT 1357.020 1710.640 1372.020 1988.560 ;
        RECT 1375.020 1710.640 1390.020 1988.560 ;
        RECT 1393.020 1710.640 1402.950 1988.560 ;
  END
END user_project_wrapper
END LIBRARY

