MACRO INVX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN INVX4 0 0 ;
 SIZE 3.12 BY 4.16 ;
 SYMMETRY X Y R90 ;
 SITE unithd ;
  PIN vdd
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.00000000 3965.00000000 3120.00000000 4355.00000000 ;
    END
  END vdd

  PIN gnd
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.00000000 -195.00000000 3120.00000000 195.00000000 ;
    END
  END gnd

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        POLYGON 405.00000000 730.00000000 405.00000000 960.00000000 450.00000000 960.00000000 450.00000000 3200.00000000 405.00000000 3200.00000000 405.00000000 3430.00000000 635.00000000 3430.00000000 635.00000000 3200.00000000 590.00000000 3200.00000000 590.00000000 960.00000000 635.00000000 960.00000000 635.00000000 915.00000000 2485.00000000 915.00000000 2485.00000000 960.00000000 2530.00000000 960.00000000 2530.00000000 3200.00000000 2485.00000000 3200.00000000 2485.00000000 3430.00000000 2715.00000000 3430.00000000 2715.00000000 3200.00000000 2670.00000000 3200.00000000 2670.00000000 960.00000000 2715.00000000 960.00000000 2715.00000000 730.00000000 2485.00000000 730.00000000 2485.00000000 775.00000000 635.00000000 775.00000000 635.00000000 730.00000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        POLYGON 925.00000000 1120.00000000 925.00000000 1350.00000000 1155.00000000 1350.00000000 1155.00000000 1305.00000000 1965.00000000 1305.00000000 1965.00000000 1350.00000000 2010.00000000 1350.00000000 2010.00000000 2810.00000000 1965.00000000 2810.00000000 1965.00000000 2855.00000000 1155.00000000 2855.00000000 1155.00000000 2810.00000000 925.00000000 2810.00000000 925.00000000 3040.00000000 1155.00000000 3040.00000000 1155.00000000 2995.00000000 1965.00000000 2995.00000000 1965.00000000 3040.00000000 2195.00000000 3040.00000000 2195.00000000 2810.00000000 2150.00000000 2810.00000000 2150.00000000 1350.00000000 2195.00000000 1350.00000000 2195.00000000 1120.00000000 1965.00000000 1120.00000000 1965.00000000 1165.00000000 1155.00000000 1165.00000000 1155.00000000 1120.00000000 ;
    END
  END A


END INVX4
