MACRO LATCH
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN LATCH 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.48000000 6.44000000 2.96000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 6.44000000 0.24000000 ;
    END
  END GND

  PIN Q
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 5.83500000 0.39500000 6.12500000 0.68500000 ;
        RECT 4.45500000 0.93500000 4.74500000 1.22500000 ;
        RECT 4.53000000 1.22500000 4.67000000 1.47500000 ;
        RECT 4.45500000 1.47500000 4.74500000 1.76500000 ;
        RECT 4.53000000 1.76500000 4.67000000 1.91000000 ;
        RECT 5.91000000 0.68500000 6.05000000 1.91000000 ;
        RECT 4.53000000 1.91000000 6.05000000 2.01500000 ;
        RECT 4.53000000 2.01500000 6.12500000 2.05000000 ;
        RECT 5.83500000 2.05000000 6.12500000 2.30500000 ;
    END
  END Q

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.61500000 0.57500000 2.90500000 0.65000000 ;
        RECT 0.85000000 0.65000000 2.90500000 0.79000000 ;
        RECT 2.61500000 0.79000000 2.90500000 0.86500000 ;
        RECT 0.85000000 0.79000000 0.99000000 0.93500000 ;
        RECT 0.77500000 0.93500000 1.06500000 1.22500000 ;
       LAYER metal2 ;
        RECT 3.53500000 1.47500000 3.82500000 1.76500000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.69500000 0.93500000 1.98500000 1.22500000 ;
    END
  END D


END LATCH
