VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NOR3X1
  CLASS CORE ;
  FOREIGN NOR3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 5.840 2.020 6.130 2.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.320 2.020 0.610 2.310 ;
        RECT 0.390 0.690 0.530 2.020 ;
        RECT 0.320 0.610 0.610 0.690 ;
        RECT 2.160 0.610 2.450 0.690 ;
        RECT 0.320 0.470 2.450 0.610 ;
        RECT 0.320 0.400 0.610 0.470 ;
        RECT 2.160 0.400 2.450 0.470 ;
    END
  END Y
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.460 1.480 4.750 1.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.700 1.480 1.990 1.770 ;
        RECT 1.770 1.230 1.910 1.480 ;
        RECT 1.700 0.940 1.990 1.230 ;
    END
  END B
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.780 1.480 1.070 1.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.780 0.940 1.070 1.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.380 1.480 5.670 1.770 ;
    END
  END C
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.620 1.690 2.910 1.770 ;
        RECT 3.540 1.690 3.830 1.770 ;
        RECT 2.620 1.550 3.830 1.690 ;
        RECT 2.620 1.480 2.910 1.550 ;
        RECT 3.540 1.480 3.830 1.550 ;
        RECT 2.690 1.230 2.830 1.480 ;
        RECT 2.620 0.940 2.910 1.230 ;
    END
  END A
END NOR3X1
END LIBRARY

