VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OAI22X1
  CLASS CORE ;
  FOREIGN OAI22X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.320 1.960 0.610 2.030 ;
        RECT 4.000 1.960 4.290 2.030 ;
        RECT 0.320 1.820 4.290 1.960 ;
        RECT 0.320 1.740 0.610 1.820 ;
        RECT 4.000 1.740 4.290 1.820 ;
        RECT 3.080 0.790 3.370 0.860 ;
        RECT 4.070 0.790 4.210 1.740 ;
        RECT 3.080 0.650 4.210 0.790 ;
        RECT 3.080 0.570 3.370 0.650 ;
    END
  END Y
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.780 1.090 1.070 1.640 ;
    END
  END B
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 3.540 1.350 3.830 1.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.620 0.440 2.910 0.730 ;
    END
  END D
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.620 1.350 2.910 1.640 ;
    END
  END C
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.700 1.090 1.990 1.640 ;
    END
  END A
END OAI22X1
END LIBRARY

