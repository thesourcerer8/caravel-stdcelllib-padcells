MACRO INV
 CLASS CORE ;
 ORIGIN 0.0 0.0 ;
 FOREIGN INV 0.0 0.0 ;
 SYMMETRY X Y R90 ;
 SITE unithd ;
  PIN vdd
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.00000000 3.96500000 2.08000000 4.35500000 ;
    END
  END vdd

  PIN gnd
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.00000000 -0.19500000 2.08000000 0.19500000 ;
    END
  END gnd

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        POLYGON 0.40500000 0.73000000 0.40500000 0.96000000 0.45000000 0.96000000 0.45000000 3.20000000 0.40500000 3.20000000 0.40500000 3.43000000 0.63500000 3.43000000 0.63500000 3.20000000 0.59000000 3.20000000 0.59000000 0.96000000 0.63500000 0.96000000 0.63500000 0.73000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        POLYGON 0.92500000 1.12000000 0.92500000 1.35000000 0.97000000 1.35000000 0.97000000 2.81000000 0.92500000 2.81000000 0.92500000 3.04000000 1.15500000 3.04000000 1.15500000 2.81000000 1.11000000 2.81000000 1.11000000 1.35000000 1.15500000 1.35000000 1.15500000 1.12000000 ;
    END
  END A


END INV
