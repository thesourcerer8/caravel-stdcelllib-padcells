MACRO XOR2X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN XOR2X1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.48000000 6.44000000 2.96000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 6.44000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 3.07500000 0.39500000 3.36500000 0.47000000 ;
        RECT 3.07500000 0.47000000 4.21000000 0.61000000 ;
        RECT 3.07500000 0.61000000 3.36500000 0.68500000 ;
        RECT 3.07500000 2.01500000 3.36500000 2.09000000 ;
        RECT 4.07000000 0.61000000 4.21000000 2.09000000 ;
        RECT 3.07500000 2.09000000 4.21000000 2.23000000 ;
        RECT 3.07500000 2.23000000 3.36500000 2.30500000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.61500000 0.57500000 2.90500000 0.65000000 ;
        RECT 0.85000000 0.65000000 2.90500000 0.79000000 ;
        RECT 2.61500000 0.79000000 2.90500000 0.86500000 ;
        RECT 0.85000000 0.79000000 0.99000000 0.93500000 ;
        RECT 0.77500000 0.93500000 1.06500000 1.22500000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.69500000 0.93500000 1.98500000 1.22500000 ;
       LAYER metal2 ;
        RECT 5.37500000 0.93500000 5.66500000 1.22500000 ;
       LAYER metal2 ;
        RECT 5.37500000 1.47500000 5.66500000 1.76500000 ;
    END
  END B


END XOR2X1
