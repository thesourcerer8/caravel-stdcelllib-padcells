MACRO HAX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN HAX1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.48000000 9.20000000 2.96000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 9.20000000 0.24000000 ;
    END
  END GND

  PIN YC
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.31500000 0.57000000 0.60500000 0.86000000 ;
        RECT 0.39000000 0.86000000 0.53000000 1.74000000 ;
        RECT 0.31500000 1.74000000 0.60500000 2.03000000 ;
    END
  END YC

  PIN YS
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 7.67500000 0.57000000 7.96500000 0.86000000 ;
    END
  END YS

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.69000000 1.03500000 5.59000000 1.09000000 ;
        RECT 2.61500000 1.09000000 5.66500000 1.17500000 ;
        RECT 2.61500000 1.17500000 2.90500000 1.64000000 ;
        RECT 5.37500000 1.17500000 5.66500000 1.64000000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 3.53500000 1.35000000 3.82500000 1.64000000 ;
       LAYER metal2 ;
        RECT 6.29500000 1.09000000 6.58500000 1.64000000 ;
       LAYER metal2 ;
        RECT 6.29500000 1.09000000 6.58500000 1.64000000 ;
    END
  END A


END HAX1
