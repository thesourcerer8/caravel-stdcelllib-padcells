MACRO BUFX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN BUFX4 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.48000000 3.68000000 2.96000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 3.68000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.15500000 0.57000000 2.44500000 0.77500000 ;
        RECT 2.15500000 0.77500000 3.29000000 0.86000000 ;
        RECT 2.23000000 0.86000000 3.29000000 0.91500000 ;
        RECT 2.15500000 1.74000000 2.44500000 1.81500000 ;
        RECT 3.15000000 0.91500000 3.29000000 1.81500000 ;
        RECT 2.15500000 1.81500000 3.29000000 1.95500000 ;
        RECT 2.15500000 1.95500000 2.44500000 2.03000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.77500000 0.96000000 1.06500000 1.25000000 ;
    END
  END A


END BUFX4
