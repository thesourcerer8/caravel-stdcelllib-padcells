MACRO NOR3X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NOR3X1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.48000000 6.44000000 2.96000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 6.44000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.31500000 0.39500000 0.60500000 0.47000000 ;
        RECT 2.15500000 0.39500000 2.44500000 0.47000000 ;
        RECT 0.31500000 0.47000000 2.44500000 0.61000000 ;
        RECT 0.31500000 0.61000000 0.60500000 0.68500000 ;
        RECT 2.15500000 0.61000000 2.44500000 0.68500000 ;
        RECT 0.39000000 0.68500000 0.53000000 2.01500000 ;
        RECT 0.31500000 2.01500000 0.60500000 2.30500000 ;
       LAYER metal2 ;
        RECT 5.83500000 2.01500000 6.12500000 2.30500000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.69500000 0.93500000 1.98500000 1.22500000 ;
        RECT 1.77000000 1.22500000 1.91000000 1.47500000 ;
        RECT 1.69500000 1.47500000 1.98500000 1.76500000 ;
       LAYER metal2 ;
        RECT 4.45500000 1.47500000 4.74500000 1.76500000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 5.37500000 1.47500000 5.66500000 1.76500000 ;
       LAYER metal2 ;
        RECT 0.77500000 0.93500000 1.06500000 1.22500000 ;
       LAYER metal2 ;
        RECT 0.77500000 1.47500000 1.06500000 1.76500000 ;
    END
  END C

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.61500000 0.93500000 2.90500000 1.22500000 ;
        RECT 2.69000000 1.22500000 2.83000000 1.47500000 ;
        RECT 2.61500000 1.47500000 2.90500000 1.55000000 ;
        RECT 3.53500000 1.47500000 3.82500000 1.55000000 ;
        RECT 2.61500000 1.55000000 3.82500000 1.69000000 ;
        RECT 2.61500000 1.69000000 2.90500000 1.76500000 ;
        RECT 3.53500000 1.69000000 3.82500000 1.76500000 ;
    END
  END A


END NOR3X1
